`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input dl_reset,
    input all_finish,
    input dl_clock);

    wire [3:0] proc_0_data_FIFO_blk;
    wire [3:0] proc_0_data_PIPO_blk;
    wire [3:0] proc_0_start_FIFO_blk;
    wire [3:0] proc_0_TLF_FIFO_blk;
    wire [3:0] proc_0_input_sync_blk;
    wire [3:0] proc_0_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_0;
    reg [3:0] proc_dep_vld_vec_0_reg;
    wire [3:0] in_chan_dep_vld_vec_0;
    wire [43:0] in_chan_dep_data_vec_0;
    wire [3:0] token_in_vec_0;
    wire [3:0] out_chan_dep_vld_vec_0;
    wire [10:0] out_chan_dep_data_0;
    wire [3:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [10:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [10:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_3_0;
    wire [10:0] dep_chan_data_3_0;
    wire token_3_0;
    wire dep_chan_vld_4_0;
    wire [10:0] dep_chan_data_4_0;
    wire token_4_0;
    wire [3:0] proc_1_data_FIFO_blk;
    wire [3:0] proc_1_data_PIPO_blk;
    wire [3:0] proc_1_start_FIFO_blk;
    wire [3:0] proc_1_TLF_FIFO_blk;
    wire [3:0] proc_1_input_sync_blk;
    wire [3:0] proc_1_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_1;
    reg [3:0] proc_dep_vld_vec_1_reg;
    wire [3:0] in_chan_dep_vld_vec_1;
    wire [43:0] in_chan_dep_data_vec_1;
    wire [3:0] token_in_vec_1;
    wire [3:0] out_chan_dep_vld_vec_1;
    wire [10:0] out_chan_dep_data_1;
    wire [3:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [10:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [10:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_3_1;
    wire [10:0] dep_chan_data_3_1;
    wire token_3_1;
    wire dep_chan_vld_5_1;
    wire [10:0] dep_chan_data_5_1;
    wire token_5_1;
    wire [3:0] proc_2_data_FIFO_blk;
    wire [3:0] proc_2_data_PIPO_blk;
    wire [3:0] proc_2_start_FIFO_blk;
    wire [3:0] proc_2_TLF_FIFO_blk;
    wire [3:0] proc_2_input_sync_blk;
    wire [3:0] proc_2_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_2;
    reg [3:0] proc_dep_vld_vec_2_reg;
    wire [3:0] in_chan_dep_vld_vec_2;
    wire [43:0] in_chan_dep_data_vec_2;
    wire [3:0] token_in_vec_2;
    wire [3:0] out_chan_dep_vld_vec_2;
    wire [10:0] out_chan_dep_data_2;
    wire [3:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [10:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [10:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [10:0] dep_chan_data_3_2;
    wire token_3_2;
    wire dep_chan_vld_4_2;
    wire [10:0] dep_chan_data_4_2;
    wire token_4_2;
    wire [3:0] proc_3_data_FIFO_blk;
    wire [3:0] proc_3_data_PIPO_blk;
    wire [3:0] proc_3_start_FIFO_blk;
    wire [3:0] proc_3_TLF_FIFO_blk;
    wire [3:0] proc_3_input_sync_blk;
    wire [3:0] proc_3_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_3;
    reg [3:0] proc_dep_vld_vec_3_reg;
    wire [3:0] in_chan_dep_vld_vec_3;
    wire [43:0] in_chan_dep_data_vec_3;
    wire [3:0] token_in_vec_3;
    wire [3:0] out_chan_dep_vld_vec_3;
    wire [10:0] out_chan_dep_data_3;
    wire [3:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_0_3;
    wire [10:0] dep_chan_data_0_3;
    wire token_0_3;
    wire dep_chan_vld_1_3;
    wire [10:0] dep_chan_data_1_3;
    wire token_1_3;
    wire dep_chan_vld_2_3;
    wire [10:0] dep_chan_data_2_3;
    wire token_2_3;
    wire dep_chan_vld_5_3;
    wire [10:0] dep_chan_data_5_3;
    wire token_5_3;
    wire [3:0] proc_4_data_FIFO_blk;
    wire [3:0] proc_4_data_PIPO_blk;
    wire [3:0] proc_4_start_FIFO_blk;
    wire [3:0] proc_4_TLF_FIFO_blk;
    wire [3:0] proc_4_input_sync_blk;
    wire [3:0] proc_4_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_4;
    reg [3:0] proc_dep_vld_vec_4_reg;
    wire [3:0] in_chan_dep_vld_vec_4;
    wire [43:0] in_chan_dep_data_vec_4;
    wire [3:0] token_in_vec_4;
    wire [3:0] out_chan_dep_vld_vec_4;
    wire [10:0] out_chan_dep_data_4;
    wire [3:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_0_4;
    wire [10:0] dep_chan_data_0_4;
    wire token_0_4;
    wire dep_chan_vld_2_4;
    wire [10:0] dep_chan_data_2_4;
    wire token_2_4;
    wire dep_chan_vld_6_4;
    wire [10:0] dep_chan_data_6_4;
    wire token_6_4;
    wire dep_chan_vld_8_4;
    wire [10:0] dep_chan_data_8_4;
    wire token_8_4;
    wire [3:0] proc_5_data_FIFO_blk;
    wire [3:0] proc_5_data_PIPO_blk;
    wire [3:0] proc_5_start_FIFO_blk;
    wire [3:0] proc_5_TLF_FIFO_blk;
    wire [3:0] proc_5_input_sync_blk;
    wire [3:0] proc_5_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_5;
    reg [3:0] proc_dep_vld_vec_5_reg;
    wire [3:0] in_chan_dep_vld_vec_5;
    wire [43:0] in_chan_dep_data_vec_5;
    wire [3:0] token_in_vec_5;
    wire [3:0] out_chan_dep_vld_vec_5;
    wire [10:0] out_chan_dep_data_5;
    wire [3:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_1_5;
    wire [10:0] dep_chan_data_1_5;
    wire token_1_5;
    wire dep_chan_vld_3_5;
    wire [10:0] dep_chan_data_3_5;
    wire token_3_5;
    wire dep_chan_vld_7_5;
    wire [10:0] dep_chan_data_7_5;
    wire token_7_5;
    wire dep_chan_vld_9_5;
    wire [10:0] dep_chan_data_9_5;
    wire token_9_5;
    wire [0:0] proc_6_data_FIFO_blk;
    wire [0:0] proc_6_data_PIPO_blk;
    wire [0:0] proc_6_start_FIFO_blk;
    wire [0:0] proc_6_TLF_FIFO_blk;
    wire [0:0] proc_6_input_sync_blk;
    wire [0:0] proc_6_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_6;
    reg [0:0] proc_dep_vld_vec_6_reg;
    wire [1:0] in_chan_dep_vld_vec_6;
    wire [21:0] in_chan_dep_data_vec_6;
    wire [1:0] token_in_vec_6;
    wire [0:0] out_chan_dep_vld_vec_6;
    wire [10:0] out_chan_dep_data_6;
    wire [0:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_4_6;
    wire [10:0] dep_chan_data_4_6;
    wire token_4_6;
    wire dep_chan_vld_8_6;
    wire [10:0] dep_chan_data_8_6;
    wire token_8_6;
    wire [0:0] proc_7_data_FIFO_blk;
    wire [0:0] proc_7_data_PIPO_blk;
    wire [0:0] proc_7_start_FIFO_blk;
    wire [0:0] proc_7_TLF_FIFO_blk;
    wire [0:0] proc_7_input_sync_blk;
    wire [0:0] proc_7_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_7;
    reg [0:0] proc_dep_vld_vec_7_reg;
    wire [1:0] in_chan_dep_vld_vec_7;
    wire [21:0] in_chan_dep_data_vec_7;
    wire [1:0] token_in_vec_7;
    wire [0:0] out_chan_dep_vld_vec_7;
    wire [10:0] out_chan_dep_data_7;
    wire [0:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_5_7;
    wire [10:0] dep_chan_data_5_7;
    wire token_5_7;
    wire dep_chan_vld_9_7;
    wire [10:0] dep_chan_data_9_7;
    wire token_9_7;
    wire [2:0] proc_8_data_FIFO_blk;
    wire [2:0] proc_8_data_PIPO_blk;
    wire [2:0] proc_8_start_FIFO_blk;
    wire [2:0] proc_8_TLF_FIFO_blk;
    wire [2:0] proc_8_input_sync_blk;
    wire [2:0] proc_8_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_8;
    reg [2:0] proc_dep_vld_vec_8_reg;
    wire [1:0] in_chan_dep_vld_vec_8;
    wire [21:0] in_chan_dep_data_vec_8;
    wire [1:0] token_in_vec_8;
    wire [2:0] out_chan_dep_vld_vec_8;
    wire [10:0] out_chan_dep_data_8;
    wire [2:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_4_8;
    wire [10:0] dep_chan_data_4_8;
    wire token_4_8;
    wire dep_chan_vld_10_8;
    wire [10:0] dep_chan_data_10_8;
    wire token_10_8;
    wire [2:0] proc_9_data_FIFO_blk;
    wire [2:0] proc_9_data_PIPO_blk;
    wire [2:0] proc_9_start_FIFO_blk;
    wire [2:0] proc_9_TLF_FIFO_blk;
    wire [2:0] proc_9_input_sync_blk;
    wire [2:0] proc_9_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_9;
    reg [2:0] proc_dep_vld_vec_9_reg;
    wire [1:0] in_chan_dep_vld_vec_9;
    wire [21:0] in_chan_dep_data_vec_9;
    wire [1:0] token_in_vec_9;
    wire [2:0] out_chan_dep_vld_vec_9;
    wire [10:0] out_chan_dep_data_9;
    wire [2:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_5_9;
    wire [10:0] dep_chan_data_5_9;
    wire token_5_9;
    wire dep_chan_vld_10_9;
    wire [10:0] dep_chan_data_10_9;
    wire token_10_9;
    wire [1:0] proc_10_data_FIFO_blk;
    wire [1:0] proc_10_data_PIPO_blk;
    wire [1:0] proc_10_start_FIFO_blk;
    wire [1:0] proc_10_TLF_FIFO_blk;
    wire [1:0] proc_10_input_sync_blk;
    wire [1:0] proc_10_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_10;
    reg [1:0] proc_dep_vld_vec_10_reg;
    wire [1:0] in_chan_dep_vld_vec_10;
    wire [21:0] in_chan_dep_data_vec_10;
    wire [1:0] token_in_vec_10;
    wire [1:0] out_chan_dep_vld_vec_10;
    wire [10:0] out_chan_dep_data_10;
    wire [1:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_8_10;
    wire [10:0] dep_chan_data_8_10;
    wire token_8_10;
    wire dep_chan_vld_9_10;
    wire [10:0] dep_chan_data_9_10;
    wire token_9_10;
    wire [10:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    wire [10:0] origin;

    reg ap_done_reg_0;// for module AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_done & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_continue;
        end
    end

    reg ap_done_reg_1;// for module AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_done & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_continue;
        end
    end

reg [15:0] trans_in_cnt_0;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_0 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.start_write == 1'b1) begin
        trans_in_cnt_0 <= trans_in_cnt_0 + 16'h1;
    end
    else begin
        trans_in_cnt_0 <= trans_in_cnt_0;
    end
end

reg [15:0] trans_out_cnt_0;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_0 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_done == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_continue == 1'b1) begin
        trans_out_cnt_0 <= trans_out_cnt_0 + 16'h1;
    end
    else begin
        trans_out_cnt_0 <= trans_out_cnt_0;
    end
end

reg [15:0] trans_in_cnt_1;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_1 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.start_write == 1'b1) begin
        trans_in_cnt_1 <= trans_in_cnt_1 + 16'h1;
    end
    else begin
        trans_in_cnt_1 <= trans_in_cnt_1;
    end
end

reg [15:0] trans_out_cnt_1;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_1 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_done == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_continue == 1'b1) begin
        trans_out_cnt_1 <= trans_out_cnt_1 + 16'h1;
    end
    else begin
        trans_out_cnt_1 <= trans_out_cnt_1;
    end
end

reg [15:0] trans_in_cnt_2;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_2 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.start_write == 1'b1) begin
        trans_in_cnt_2 <= trans_in_cnt_2 + 16'h1;
    end
    else begin
        trans_in_cnt_2 <= trans_in_cnt_2;
    end
end

reg [15:0] trans_out_cnt_2;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_2 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_done == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_continue == 1'b1) begin
        trans_out_cnt_2 <= trans_out_cnt_2 + 16'h1;
    end
    else begin
        trans_out_cnt_2 <= trans_out_cnt_2;
    end
end

reg [15:0] trans_in_cnt_3;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_3 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.start_write == 1'b1) begin
        trans_in_cnt_3 <= trans_in_cnt_3 + 16'h1;
    end
    else begin
        trans_in_cnt_3 <= trans_in_cnt_3;
    end
end

reg [15:0] trans_out_cnt_3;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_3 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.ap_done == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.ap_continue == 1'b1) begin
        trans_out_cnt_3 <= trans_out_cnt_3 + 16'h1;
    end
    else begin
        trans_out_cnt_3 <= trans_out_cnt_3;
    end
end

reg [15:0] trans_in_cnt_4;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_4 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.start_write == 1'b1) begin
        trans_in_cnt_4 <= trans_in_cnt_4 + 16'h1;
    end
    else begin
        trans_in_cnt_4 <= trans_in_cnt_4;
    end
end

reg [15:0] trans_out_cnt_4;// for process AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_4 <= 16'h0;
    end
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_done == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_continue == 1'b1) begin
        trans_out_cnt_4 <= trans_out_cnt_4 + 16'h1;
    end
    else begin
        trans_out_cnt_4 <= trans_out_cnt_4;
    end
end

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
    AESL_deadlock_detect_unit #(11, 0, 4, 4) AESL_deadlock_detect_unit_0 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_3_blk_n);
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0;
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    assign proc_0_data_FIFO_blk[1] = 1'b0;
    assign proc_0_data_PIPO_blk[1] = 1'b0;
    assign proc_0_start_FIFO_blk[1] = 1'b0;
    assign proc_0_TLF_FIFO_blk[1] = 1'b0;
    assign proc_0_input_sync_blk[1] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready);
    assign proc_0_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (proc_0_data_FIFO_blk[1] | proc_0_data_PIPO_blk[1] | proc_0_start_FIFO_blk[1] | proc_0_TLF_FIFO_blk[1] | proc_0_input_sync_blk[1] | proc_0_output_sync_blk[1]);
    assign proc_0_data_FIFO_blk[2] = 1'b0;
    assign proc_0_data_PIPO_blk[2] = 1'b0;
    assign proc_0_start_FIFO_blk[2] = 1'b0;
    assign proc_0_TLF_FIFO_blk[2] = 1'b0;
    assign proc_0_input_sync_blk[2] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready);
    assign proc_0_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (proc_0_data_FIFO_blk[2] | proc_0_data_PIPO_blk[2] | proc_0_start_FIFO_blk[2] | proc_0_TLF_FIFO_blk[2] | proc_0_input_sync_blk[2] | proc_0_output_sync_blk[2]);
    assign proc_0_data_FIFO_blk[3] = 1'b0;
    assign proc_0_data_PIPO_blk[3] = 1'b0;
    assign proc_0_start_FIFO_blk[3] = 1'b0;
    assign proc_0_TLF_FIFO_blk[3] = 1'b0;
    assign proc_0_input_sync_blk[3] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready);
    assign proc_0_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_0[3] = dl_detect_out ? proc_dep_vld_vec_0_reg[3] : (proc_0_data_FIFO_blk[3] | proc_0_data_PIPO_blk[3] | proc_0_start_FIFO_blk[3] | proc_0_TLF_FIFO_blk[3] | proc_0_input_sync_blk[3] | proc_0_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[10 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[21 : 11] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_3_0;
    assign in_chan_dep_data_vec_0[32 : 22] = dep_chan_data_3_0;
    assign token_in_vec_0[2] = token_3_0;
    assign in_chan_dep_vld_vec_0[3] = dep_chan_vld_4_0;
    assign in_chan_dep_data_vec_0[43 : 33] = dep_chan_data_4_0;
    assign token_in_vec_0[3] = token_4_0;
    assign dep_chan_vld_0_4 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_4 = out_chan_dep_data_0;
    assign token_0_4 = token_out_vec_0[0];
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[1];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[2];
    assign dep_chan_vld_0_3 = out_chan_dep_vld_vec_0[3];
    assign dep_chan_data_0_3 = out_chan_dep_data_0;
    assign token_0_3 = token_out_vec_0[3];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0
    AESL_deadlock_detect_unit #(11, 1, 4, 4) AESL_deadlock_detect_unit_1 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_3_blk_n);
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_read);
    assign proc_1_TLF_FIFO_blk[0] = 1'b0;
    assign proc_1_input_sync_blk[0] = 1'b0;
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    assign proc_1_data_FIFO_blk[1] = 1'b0;
    assign proc_1_data_PIPO_blk[1] = 1'b0;
    assign proc_1_start_FIFO_blk[1] = 1'b0;
    assign proc_1_TLF_FIFO_blk[1] = 1'b0;
    assign proc_1_input_sync_blk[1] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready);
    assign proc_1_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (proc_1_data_FIFO_blk[1] | proc_1_data_PIPO_blk[1] | proc_1_start_FIFO_blk[1] | proc_1_TLF_FIFO_blk[1] | proc_1_input_sync_blk[1] | proc_1_output_sync_blk[1]);
    assign proc_1_data_FIFO_blk[2] = 1'b0;
    assign proc_1_data_PIPO_blk[2] = 1'b0;
    assign proc_1_start_FIFO_blk[2] = 1'b0;
    assign proc_1_TLF_FIFO_blk[2] = 1'b0;
    assign proc_1_input_sync_blk[2] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready);
    assign proc_1_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (proc_1_data_FIFO_blk[2] | proc_1_data_PIPO_blk[2] | proc_1_start_FIFO_blk[2] | proc_1_TLF_FIFO_blk[2] | proc_1_input_sync_blk[2] | proc_1_output_sync_blk[2]);
    assign proc_1_data_FIFO_blk[3] = 1'b0;
    assign proc_1_data_PIPO_blk[3] = 1'b0;
    assign proc_1_start_FIFO_blk[3] = 1'b0;
    assign proc_1_TLF_FIFO_blk[3] = 1'b0;
    assign proc_1_input_sync_blk[3] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready);
    assign proc_1_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (proc_1_data_FIFO_blk[3] | proc_1_data_PIPO_blk[3] | proc_1_start_FIFO_blk[3] | proc_1_TLF_FIFO_blk[3] | proc_1_input_sync_blk[3] | proc_1_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[10 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[21 : 11] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_3_1;
    assign in_chan_dep_data_vec_1[32 : 22] = dep_chan_data_3_1;
    assign token_in_vec_1[2] = token_3_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_5_1;
    assign in_chan_dep_data_vec_1[43 : 33] = dep_chan_data_5_1;
    assign token_in_vec_1[3] = token_5_1;
    assign dep_chan_vld_1_5 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_5 = out_chan_dep_data_1;
    assign token_1_5 = token_out_vec_1[0];
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[1];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[2];
    assign dep_chan_vld_1_3 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_3 = out_chan_dep_data_1;
    assign token_1_3 = token_out_vec_1[3];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0
    AESL_deadlock_detect_unit #(11, 2, 4, 4) AESL_deadlock_detect_unit_2 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_2_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_3_blk_n);
    assign proc_2_data_PIPO_blk[0] = 1'b0;
    assign proc_2_start_FIFO_blk[0] = 1'b0;
    assign proc_2_TLF_FIFO_blk[0] = 1'b0;
    assign proc_2_input_sync_blk[0] = 1'b0;
    assign proc_2_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (proc_2_data_FIFO_blk[0] | proc_2_data_PIPO_blk[0] | proc_2_start_FIFO_blk[0] | proc_2_TLF_FIFO_blk[0] | proc_2_input_sync_blk[0] | proc_2_output_sync_blk[0]);
    assign proc_2_data_FIFO_blk[1] = 1'b0;
    assign proc_2_data_PIPO_blk[1] = 1'b0;
    assign proc_2_start_FIFO_blk[1] = 1'b0;
    assign proc_2_TLF_FIFO_blk[1] = 1'b0;
    assign proc_2_input_sync_blk[1] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready);
    assign proc_2_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (proc_2_data_FIFO_blk[1] | proc_2_data_PIPO_blk[1] | proc_2_start_FIFO_blk[1] | proc_2_TLF_FIFO_blk[1] | proc_2_input_sync_blk[1] | proc_2_output_sync_blk[1]);
    assign proc_2_data_FIFO_blk[2] = 1'b0;
    assign proc_2_data_PIPO_blk[2] = 1'b0;
    assign proc_2_start_FIFO_blk[2] = 1'b0;
    assign proc_2_TLF_FIFO_blk[2] = 1'b0;
    assign proc_2_input_sync_blk[2] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready);
    assign proc_2_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (proc_2_data_FIFO_blk[2] | proc_2_data_PIPO_blk[2] | proc_2_start_FIFO_blk[2] | proc_2_TLF_FIFO_blk[2] | proc_2_input_sync_blk[2] | proc_2_output_sync_blk[2]);
    assign proc_2_data_FIFO_blk[3] = 1'b0;
    assign proc_2_data_PIPO_blk[3] = 1'b0;
    assign proc_2_start_FIFO_blk[3] = 1'b0;
    assign proc_2_TLF_FIFO_blk[3] = 1'b0;
    assign proc_2_input_sync_blk[3] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready);
    assign proc_2_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_2[3] = dl_detect_out ? proc_dep_vld_vec_2_reg[3] : (proc_2_data_FIFO_blk[3] | proc_2_data_PIPO_blk[3] | proc_2_start_FIFO_blk[3] | proc_2_TLF_FIFO_blk[3] | proc_2_input_sync_blk[3] | proc_2_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[10 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[21 : 11] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[32 : 22] = dep_chan_data_3_2;
    assign token_in_vec_2[2] = token_3_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_4_2;
    assign in_chan_dep_data_vec_2[43 : 33] = dep_chan_data_4_2;
    assign token_in_vec_2[3] = token_4_2;
    assign dep_chan_vld_2_4 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_4 = out_chan_dep_data_2;
    assign token_2_4 = token_out_vec_2[0];
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[1];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[2];
    assign dep_chan_vld_2_3 = out_chan_dep_vld_vec_2[3];
    assign dep_chan_data_2_3 = out_chan_dep_data_2;
    assign token_2_3 = token_out_vec_2[3];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0
    AESL_deadlock_detect_unit #(11, 3, 4, 4) AESL_deadlock_detect_unit_3 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_3_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_3_blk_n);
    assign proc_3_data_PIPO_blk[0] = 1'b0;
    assign proc_3_start_FIFO_blk[0] = 1'b0;
    assign proc_3_TLF_FIFO_blk[0] = 1'b0;
    assign proc_3_input_sync_blk[0] = 1'b0;
    assign proc_3_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (proc_3_data_FIFO_blk[0] | proc_3_data_PIPO_blk[0] | proc_3_start_FIFO_blk[0] | proc_3_TLF_FIFO_blk[0] | proc_3_input_sync_blk[0] | proc_3_output_sync_blk[0]);
    assign proc_3_data_FIFO_blk[1] = 1'b0;
    assign proc_3_data_PIPO_blk[1] = 1'b0;
    assign proc_3_start_FIFO_blk[1] = 1'b0;
    assign proc_3_TLF_FIFO_blk[1] = 1'b0;
    assign proc_3_input_sync_blk[1] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready);
    assign proc_3_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (proc_3_data_FIFO_blk[1] | proc_3_data_PIPO_blk[1] | proc_3_start_FIFO_blk[1] | proc_3_TLF_FIFO_blk[1] | proc_3_input_sync_blk[1] | proc_3_output_sync_blk[1]);
    assign proc_3_data_FIFO_blk[2] = 1'b0;
    assign proc_3_data_PIPO_blk[2] = 1'b0;
    assign proc_3_start_FIFO_blk[2] = 1'b0;
    assign proc_3_TLF_FIFO_blk[2] = 1'b0;
    assign proc_3_input_sync_blk[2] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready);
    assign proc_3_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (proc_3_data_FIFO_blk[2] | proc_3_data_PIPO_blk[2] | proc_3_start_FIFO_blk[2] | proc_3_TLF_FIFO_blk[2] | proc_3_input_sync_blk[2] | proc_3_output_sync_blk[2]);
    assign proc_3_data_FIFO_blk[3] = 1'b0;
    assign proc_3_data_PIPO_blk[3] = 1'b0;
    assign proc_3_start_FIFO_blk[3] = 1'b0;
    assign proc_3_TLF_FIFO_blk[3] = 1'b0;
    assign proc_3_input_sync_blk[3] = 1'b0 | (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready);
    assign proc_3_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_3[3] = dl_detect_out ? proc_dep_vld_vec_3_reg[3] : (proc_3_data_FIFO_blk[3] | proc_3_data_PIPO_blk[3] | proc_3_start_FIFO_blk[3] | proc_3_TLF_FIFO_blk[3] | proc_3_input_sync_blk[3] | proc_3_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_0_3;
    assign in_chan_dep_data_vec_3[10 : 0] = dep_chan_data_0_3;
    assign token_in_vec_3[0] = token_0_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_1_3;
    assign in_chan_dep_data_vec_3[21 : 11] = dep_chan_data_1_3;
    assign token_in_vec_3[1] = token_1_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_2_3;
    assign in_chan_dep_data_vec_3[32 : 22] = dep_chan_data_2_3;
    assign token_in_vec_3[2] = token_2_3;
    assign in_chan_dep_vld_vec_3[3] = dep_chan_vld_5_3;
    assign in_chan_dep_data_vec_3[43 : 33] = dep_chan_data_5_3;
    assign token_in_vec_3[3] = token_5_3;
    assign dep_chan_vld_3_5 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_5 = out_chan_dep_data_3;
    assign token_3_5 = token_out_vec_3[0];
    assign dep_chan_vld_3_0 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_0 = out_chan_dep_data_3;
    assign token_3_0 = token_out_vec_3[1];
    assign dep_chan_vld_3_1 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_1 = out_chan_dep_data_3;
    assign token_3_1 = token_out_vec_3[2];
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[3];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[3];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
    AESL_deadlock_detect_unit #(11, 4, 4, 4) AESL_deadlock_detect_unit_4 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_4_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_3_blk_n);
    assign proc_4_data_PIPO_blk[0] = 1'b0;
    assign proc_4_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_write);
    assign proc_4_TLF_FIFO_blk[0] = 1'b0;
    assign proc_4_input_sync_blk[0] = 1'b0;
    assign proc_4_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (proc_4_data_FIFO_blk[0] | proc_4_data_PIPO_blk[0] | proc_4_start_FIFO_blk[0] | proc_4_TLF_FIFO_blk[0] | proc_4_input_sync_blk[0] | proc_4_output_sync_blk[0]);
    assign proc_4_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_value_0_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_value_0_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_value_0_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_value_0_3_blk_n);
    assign proc_4_data_PIPO_blk[1] = 1'b0;
    assign proc_4_start_FIFO_blk[1] = 1'b0;
    assign proc_4_TLF_FIFO_blk[1] = 1'b0;
    assign proc_4_input_sync_blk[1] = 1'b0;
    assign proc_4_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (proc_4_data_FIFO_blk[1] | proc_4_data_PIPO_blk[1] | proc_4_start_FIFO_blk[1] | proc_4_TLF_FIFO_blk[1] | proc_4_input_sync_blk[1] | proc_4_output_sync_blk[1]);
    assign proc_4_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.k_proj_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.q_proj_0_blk_n);
    assign proc_4_data_PIPO_blk[2] = 1'b0;
    assign proc_4_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_read);
    assign proc_4_TLF_FIFO_blk[2] = 1'b0;
    assign proc_4_input_sync_blk[2] = 1'b0;
    assign proc_4_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_4[2] = dl_detect_out ? proc_dep_vld_vec_4_reg[2] : (proc_4_data_FIFO_blk[2] | proc_4_data_PIPO_blk[2] | proc_4_start_FIFO_blk[2] | proc_4_TLF_FIFO_blk[2] | proc_4_input_sync_blk[2] | proc_4_output_sync_blk[2]);
    assign proc_4_data_FIFO_blk[3] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.v_proj_0_blk_n);
    assign proc_4_data_PIPO_blk[3] = 1'b0;
    assign proc_4_start_FIFO_blk[3] = 1'b0;
    assign proc_4_TLF_FIFO_blk[3] = 1'b0;
    assign proc_4_input_sync_blk[3] = 1'b0;
    assign proc_4_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_4[3] = dl_detect_out ? proc_dep_vld_vec_4_reg[3] : (proc_4_data_FIFO_blk[3] | proc_4_data_PIPO_blk[3] | proc_4_start_FIFO_blk[3] | proc_4_TLF_FIFO_blk[3] | proc_4_input_sync_blk[3] | proc_4_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_0_4;
    assign in_chan_dep_data_vec_4[10 : 0] = dep_chan_data_0_4;
    assign token_in_vec_4[0] = token_0_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_2_4;
    assign in_chan_dep_data_vec_4[21 : 11] = dep_chan_data_2_4;
    assign token_in_vec_4[1] = token_2_4;
    assign in_chan_dep_vld_vec_4[2] = dep_chan_vld_6_4;
    assign in_chan_dep_data_vec_4[32 : 22] = dep_chan_data_6_4;
    assign token_in_vec_4[2] = token_6_4;
    assign in_chan_dep_vld_vec_4[3] = dep_chan_vld_8_4;
    assign in_chan_dep_data_vec_4[43 : 33] = dep_chan_data_8_4;
    assign token_in_vec_4[3] = token_8_4;
    assign dep_chan_vld_4_0 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_0 = out_chan_dep_data_4;
    assign token_4_0 = token_out_vec_4[0];
    assign dep_chan_vld_4_2 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_2 = out_chan_dep_data_4;
    assign token_4_2 = token_out_vec_4[1];
    assign dep_chan_vld_4_6 = out_chan_dep_vld_vec_4[2];
    assign dep_chan_data_4_6 = out_chan_dep_data_4;
    assign token_4_6 = token_out_vec_4[2];
    assign dep_chan_vld_4_8 = out_chan_dep_vld_vec_4[3];
    assign dep_chan_data_4_8 = out_chan_dep_data_4;
    assign token_4_8 = token_out_vec_4[3];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0
    AESL_deadlock_detect_unit #(11, 5, 4, 4) AESL_deadlock_detect_unit_5 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_5_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_query_1_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_query_1_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_query_1_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_query_1_3_blk_n);
    assign proc_5_data_PIPO_blk[0] = 1'b0;
    assign proc_5_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_write);
    assign proc_5_TLF_FIFO_blk[0] = 1'b0;
    assign proc_5_input_sync_blk[0] = 1'b0;
    assign proc_5_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (proc_5_data_FIFO_blk[0] | proc_5_data_PIPO_blk[0] | proc_5_start_FIFO_blk[0] | proc_5_TLF_FIFO_blk[0] | proc_5_input_sync_blk[0] | proc_5_output_sync_blk[0]);
    assign proc_5_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_value_1_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_value_1_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_value_1_2_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_value_1_3_blk_n);
    assign proc_5_data_PIPO_blk[1] = 1'b0;
    assign proc_5_start_FIFO_blk[1] = 1'b0;
    assign proc_5_TLF_FIFO_blk[1] = 1'b0;
    assign proc_5_input_sync_blk[1] = 1'b0;
    assign proc_5_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (proc_5_data_FIFO_blk[1] | proc_5_data_PIPO_blk[1] | proc_5_start_FIFO_blk[1] | proc_5_TLF_FIFO_blk[1] | proc_5_input_sync_blk[1] | proc_5_output_sync_blk[1]);
    assign proc_5_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.k_proj_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.q_proj_1_blk_n);
    assign proc_5_data_PIPO_blk[2] = 1'b0;
    assign proc_5_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_read);
    assign proc_5_TLF_FIFO_blk[2] = 1'b0;
    assign proc_5_input_sync_blk[2] = 1'b0;
    assign proc_5_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (proc_5_data_FIFO_blk[2] | proc_5_data_PIPO_blk[2] | proc_5_start_FIFO_blk[2] | proc_5_TLF_FIFO_blk[2] | proc_5_input_sync_blk[2] | proc_5_output_sync_blk[2]);
    assign proc_5_data_FIFO_blk[3] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.v_proj_1_blk_n);
    assign proc_5_data_PIPO_blk[3] = 1'b0;
    assign proc_5_start_FIFO_blk[3] = 1'b0;
    assign proc_5_TLF_FIFO_blk[3] = 1'b0;
    assign proc_5_input_sync_blk[3] = 1'b0;
    assign proc_5_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_5[3] = dl_detect_out ? proc_dep_vld_vec_5_reg[3] : (proc_5_data_FIFO_blk[3] | proc_5_data_PIPO_blk[3] | proc_5_start_FIFO_blk[3] | proc_5_TLF_FIFO_blk[3] | proc_5_input_sync_blk[3] | proc_5_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_1_5;
    assign in_chan_dep_data_vec_5[10 : 0] = dep_chan_data_1_5;
    assign token_in_vec_5[0] = token_1_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_3_5;
    assign in_chan_dep_data_vec_5[21 : 11] = dep_chan_data_3_5;
    assign token_in_vec_5[1] = token_3_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_7_5;
    assign in_chan_dep_data_vec_5[32 : 22] = dep_chan_data_7_5;
    assign token_in_vec_5[2] = token_7_5;
    assign in_chan_dep_vld_vec_5[3] = dep_chan_vld_9_5;
    assign in_chan_dep_data_vec_5[43 : 33] = dep_chan_data_9_5;
    assign token_in_vec_5[3] = token_9_5;
    assign dep_chan_vld_5_1 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_1 = out_chan_dep_data_5;
    assign token_5_1 = token_out_vec_5[0];
    assign dep_chan_vld_5_3 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_3 = out_chan_dep_data_5;
    assign token_5_3 = token_out_vec_5[1];
    assign dep_chan_vld_5_7 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_7 = out_chan_dep_data_5;
    assign token_5_7 = token_out_vec_5[2];
    assign dep_chan_vld_5_9 = out_chan_dep_vld_vec_5[3];
    assign dep_chan_data_5_9 = out_chan_dep_data_5;
    assign token_5_9 = token_out_vec_5[3];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0
    AESL_deadlock_detect_unit #(11, 6, 2, 1) AESL_deadlock_detect_unit_6 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_6_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0.q_proj_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0.k_proj_0_blk_n);
    assign proc_6_data_PIPO_blk[0] = 1'b0;
    assign proc_6_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_write);
    assign proc_6_TLF_FIFO_blk[0] = 1'b0;
    assign proc_6_input_sync_blk[0] = 1'b0;
    assign proc_6_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (proc_6_data_FIFO_blk[0] | proc_6_data_PIPO_blk[0] | proc_6_start_FIFO_blk[0] | proc_6_TLF_FIFO_blk[0] | proc_6_input_sync_blk[0] | proc_6_output_sync_blk[0]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_4_6;
    assign in_chan_dep_data_vec_6[10 : 0] = dep_chan_data_4_6;
    assign token_in_vec_6[0] = token_4_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_8_6;
    assign in_chan_dep_data_vec_6[21 : 11] = dep_chan_data_8_6;
    assign token_in_vec_6[1] = token_8_6;
    assign dep_chan_vld_6_4 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_4 = out_chan_dep_data_6;
    assign token_6_4 = token_out_vec_6[0];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0
    AESL_deadlock_detect_unit #(11, 7, 2, 1) AESL_deadlock_detect_unit_7 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_7_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0.q_proj_1_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0.k_proj_1_blk_n);
    assign proc_7_data_PIPO_blk[0] = 1'b0;
    assign proc_7_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_write);
    assign proc_7_TLF_FIFO_blk[0] = 1'b0;
    assign proc_7_input_sync_blk[0] = 1'b0;
    assign proc_7_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (proc_7_data_FIFO_blk[0] | proc_7_data_PIPO_blk[0] | proc_7_start_FIFO_blk[0] | proc_7_TLF_FIFO_blk[0] | proc_7_input_sync_blk[0] | proc_7_output_sync_blk[0]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_5_7;
    assign in_chan_dep_data_vec_7[10 : 0] = dep_chan_data_5_7;
    assign token_in_vec_7[0] = token_5_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_9_7;
    assign in_chan_dep_data_vec_7[21 : 11] = dep_chan_data_9_7;
    assign token_in_vec_7[1] = token_9_7;
    assign dep_chan_vld_7_5 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_5 = out_chan_dep_data_7;
    assign token_7_5 = token_out_vec_7[0];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
    AESL_deadlock_detect_unit #(11, 8, 2, 3) AESL_deadlock_detect_unit_8 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_8_data_FIFO_blk[0] = 1'b0;
    assign proc_8_data_PIPO_blk[0] = 1'b0;
    assign proc_8_start_FIFO_blk[0] = 1'b0;
    assign proc_8_TLF_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U.if_write);
    assign proc_8_input_sync_blk[0] = 1'b0;
    assign proc_8_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (proc_8_data_FIFO_blk[0] | proc_8_data_PIPO_blk[0] | proc_8_start_FIFO_blk[0] | proc_8_TLF_FIFO_blk[0] | proc_8_input_sync_blk[0] | proc_8_output_sync_blk[0]);
    assign proc_8_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.v_proj_0_blk_n);
    assign proc_8_data_PIPO_blk[1] = 1'b0;
    assign proc_8_start_FIFO_blk[1] = 1'b0;
    assign proc_8_TLF_FIFO_blk[1] = 1'b0;
    assign proc_8_input_sync_blk[1] = 1'b0;
    assign proc_8_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (proc_8_data_FIFO_blk[1] | proc_8_data_PIPO_blk[1] | proc_8_start_FIFO_blk[1] | proc_8_TLF_FIFO_blk[1] | proc_8_input_sync_blk[1] | proc_8_output_sync_blk[1]);
    assign proc_8_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_1_blk_n);
    assign proc_8_data_PIPO_blk[2] = 1'b0;
    assign proc_8_start_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_read);
    assign proc_8_TLF_FIFO_blk[2] = 1'b0;
    assign proc_8_input_sync_blk[2] = 1'b0;
    assign proc_8_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_8[2] = dl_detect_out ? proc_dep_vld_vec_8_reg[2] : (proc_8_data_FIFO_blk[2] | proc_8_data_PIPO_blk[2] | proc_8_start_FIFO_blk[2] | proc_8_TLF_FIFO_blk[2] | proc_8_input_sync_blk[2] | proc_8_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_4_8;
    assign in_chan_dep_data_vec_8[10 : 0] = dep_chan_data_4_8;
    assign token_in_vec_8[0] = token_4_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_10_8;
    assign in_chan_dep_data_vec_8[21 : 11] = dep_chan_data_10_8;
    assign token_in_vec_8[1] = token_10_8;
    assign dep_chan_vld_8_6 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_6 = out_chan_dep_data_8;
    assign token_8_6 = token_out_vec_8[0];
    assign dep_chan_vld_8_4 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_4 = out_chan_dep_data_8;
    assign token_8_4 = token_out_vec_8[1];
    assign dep_chan_vld_8_10 = out_chan_dep_vld_vec_8[2];
    assign dep_chan_data_8_10 = out_chan_dep_data_8;
    assign token_8_10 = token_out_vec_8[2];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0
    AESL_deadlock_detect_unit #(11, 9, 2, 3) AESL_deadlock_detect_unit_9 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_9_data_FIFO_blk[0] = 1'b0;
    assign proc_9_data_PIPO_blk[0] = 1'b0;
    assign proc_9_start_FIFO_blk[0] = 1'b0;
    assign proc_9_TLF_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U.if_write) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U.if_write);
    assign proc_9_input_sync_blk[0] = 1'b0;
    assign proc_9_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (proc_9_data_FIFO_blk[0] | proc_9_data_PIPO_blk[0] | proc_9_start_FIFO_blk[0] | proc_9_TLF_FIFO_blk[0] | proc_9_input_sync_blk[0] | proc_9_output_sync_blk[0]);
    assign proc_9_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.v_proj_1_blk_n);
    assign proc_9_data_PIPO_blk[1] = 1'b0;
    assign proc_9_start_FIFO_blk[1] = 1'b0;
    assign proc_9_TLF_FIFO_blk[1] = 1'b0;
    assign proc_9_input_sync_blk[1] = 1'b0;
    assign proc_9_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (proc_9_data_FIFO_blk[1] | proc_9_data_PIPO_blk[1] | proc_9_start_FIFO_blk[1] | proc_9_TLF_FIFO_blk[1] | proc_9_input_sync_blk[1] | proc_9_output_sync_blk[1]);
    assign proc_9_data_FIFO_blk[2] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.matr_out_1_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.matr_out_1_1_blk_n);
    assign proc_9_data_PIPO_blk[2] = 1'b0;
    assign proc_9_start_FIFO_blk[2] = 1'b0;
    assign proc_9_TLF_FIFO_blk[2] = 1'b0;
    assign proc_9_input_sync_blk[2] = 1'b0;
    assign proc_9_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (proc_9_data_FIFO_blk[2] | proc_9_data_PIPO_blk[2] | proc_9_start_FIFO_blk[2] | proc_9_TLF_FIFO_blk[2] | proc_9_input_sync_blk[2] | proc_9_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_5_9;
    assign in_chan_dep_data_vec_9[10 : 0] = dep_chan_data_5_9;
    assign token_in_vec_9[0] = token_5_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[21 : 11] = dep_chan_data_10_9;
    assign token_in_vec_9[1] = token_10_9;
    assign dep_chan_vld_9_7 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_7 = out_chan_dep_data_9;
    assign token_9_7 = token_out_vec_9[0];
    assign dep_chan_vld_9_5 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_5 = out_chan_dep_data_9;
    assign token_9_5 = token_out_vec_9[1];
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[2];

    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
    AESL_deadlock_detect_unit #(11, 10, 2, 2) AESL_deadlock_detect_unit_10 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_10_data_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_1_blk_n);
    assign proc_10_data_PIPO_blk[0] = 1'b0;
    assign proc_10_start_FIFO_blk[0] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_write);
    assign proc_10_TLF_FIFO_blk[0] = 1'b0;
    assign proc_10_input_sync_blk[0] = 1'b0;
    assign proc_10_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (proc_10_data_FIFO_blk[0] | proc_10_data_PIPO_blk[0] | proc_10_start_FIFO_blk[0] | proc_10_TLF_FIFO_blk[0] | proc_10_input_sync_blk[0] | proc_10_output_sync_blk[0]);
    assign proc_10_data_FIFO_blk[1] = 1'b0 | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_1_0_blk_n) | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_1_1_blk_n);
    assign proc_10_data_PIPO_blk[1] = 1'b0;
    assign proc_10_start_FIFO_blk[1] = 1'b0;
    assign proc_10_TLF_FIFO_blk[1] = 1'b0;
    assign proc_10_input_sync_blk[1] = 1'b0;
    assign proc_10_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (proc_10_data_FIFO_blk[1] | proc_10_data_PIPO_blk[1] | proc_10_start_FIFO_blk[1] | proc_10_TLF_FIFO_blk[1] | proc_10_input_sync_blk[1] | proc_10_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_8_10;
    assign in_chan_dep_data_vec_10[10 : 0] = dep_chan_data_8_10;
    assign token_in_vec_10[0] = token_8_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[21 : 11] = dep_chan_data_9_10;
    assign token_in_vec_10[1] = token_9_10;
    assign dep_chan_vld_10_8 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_8 = out_chan_dep_data_10;
    assign token_10_8 = token_out_vec_10[0];
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[1];


    wire [10:0] dl_in_vec_comb = dl_in_vec & ~{10{all_finish}};
    AESL_deadlock_report_unit #(11) AESL_deadlock_report_unit_inst (
        .dl_reset(dl_reset),
        .dl_clock(dl_clock),
        .dl_in_vec(dl_in_vec_comb),
        .trans_in_cnt_0(trans_in_cnt_0),
        .trans_out_cnt_0(trans_out_cnt_0),
        .trans_in_cnt_1(trans_in_cnt_1),
        .trans_out_cnt_1(trans_out_cnt_1),
        .trans_in_cnt_2(trans_in_cnt_2),
        .trans_out_cnt_2(trans_out_cnt_2),
        .trans_in_cnt_3(trans_in_cnt_3),
        .trans_out_cnt_3(trans_out_cnt_3),
        .trans_in_cnt_4(trans_in_cnt_4),
        .trans_out_cnt_4(trans_out_cnt_4),
        .ap_done_reg_0(ap_done_reg_0),
        .ap_done_reg_1(ap_done_reg_1),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
