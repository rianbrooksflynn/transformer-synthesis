`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input dl_reset,
    input dl_clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    input [15:0] trans_in_cnt_0,
    input [15:0] trans_out_cnt_0,
    input [15:0] trans_in_cnt_1,
    input [15:0] trans_out_cnt_1,
    input [15:0] trans_in_cnt_2,
    input [15:0] trans_out_cnt_2,
    input [15:0] trans_in_cnt_3,
    input [15:0] trans_out_cnt_3,
    input [15:0] trans_in_cnt_4,
    input [15:0] trans_out_cnt_4,
    input ap_done_reg_0,
    input ap_done_reg_1,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 3'b000;
    localparam ST_FILTER_FAKE = 3'b001;
    localparam ST_DL_DETECTED = 3'b010;
    localparam ST_DL_REPORT = 3'b100;

    reg find_df_deadlock;
    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [1352:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0";
                end
                1 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0";
                end
                2 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0";
                end
                3 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0";
                end
                4 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0";
                end
                5 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0";
                end
                6 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0";
                end
                7 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0";
                end
                8 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0";
                end
                9 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0";
                end
                10 : begin
                    proc_path = "myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [1352:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [1352:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [1448:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_3_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0',");
                        end
                    end
                    1: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.d_query_1_3_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0',");
                        end
                    end
                    0: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.d_value_0_3_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                        end
                    end
                    1: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                        end
                    end
                    3: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.d_value_1_3_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                        end
                    end
                    1: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                        end
                    end
                    2: begin
                        if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0_ap_ready & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.ap_sync_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    0: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_query_0_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0',");
                        end
                    end
                    2: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_value_0_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.d_value_0_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.k_proj_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.q_proj_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0',");
                        end
                    end
                    8: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.v_proj_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    1: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_query_1_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_query_1_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_query_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_6_U0',");
                        end
                    end
                    3: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_value_1_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.d_value_1_2_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.d_value_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    7: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.k_proj_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.q_proj_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0',");
                        end
                    end
                    9: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0.v_proj_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0.q_proj_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0.k_proj_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0',");
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0.q_proj_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.q_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0.k_proj_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.k_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0',");
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    6: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    4: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.v_proj_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_start & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0',");
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_0_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_1_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_2_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_3_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_4_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_5_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_6_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_7_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_8_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_9_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_10_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_11_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_12_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_13_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_14_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_15_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_16_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_17_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_18_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U.if_write) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.qk_mul_19_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.v_proj_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.v_proj_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.matr_out_1_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0.matr_out_1_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_0_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0',");
                        end
                    end
                    9: begin
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_1_0_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.matr_out_1_1_blk_n) begin
                            if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U' written by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U' read by process 'myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_206.matr_out_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
