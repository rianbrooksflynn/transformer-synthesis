`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [3:0] proc_dep_vld_vec_0;
    reg [3:0] proc_dep_vld_vec_0_reg;
    wire [3:0] in_chan_dep_vld_vec_0;
    wire [47:0] in_chan_dep_data_vec_0;
    wire [3:0] token_in_vec_0;
    wire [3:0] out_chan_dep_vld_vec_0;
    wire [11:0] out_chan_dep_data_0;
    wire [3:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [11:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [11:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_3_0;
    wire [11:0] dep_chan_data_3_0;
    wire token_3_0;
    wire dep_chan_vld_4_0;
    wire [11:0] dep_chan_data_4_0;
    wire token_4_0;
    wire [1:0] proc_dep_vld_vec_1;
    reg [1:0] proc_dep_vld_vec_1_reg;
    wire [1:0] in_chan_dep_vld_vec_1;
    wire [23:0] in_chan_dep_data_vec_1;
    wire [1:0] token_in_vec_1;
    wire [1:0] out_chan_dep_vld_vec_1;
    wire [11:0] out_chan_dep_data_1;
    wire [1:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [11:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_5_1;
    wire [11:0] dep_chan_data_5_1;
    wire token_5_1;
    wire [1:0] proc_dep_vld_vec_2;
    reg [1:0] proc_dep_vld_vec_2_reg;
    wire [1:0] in_chan_dep_vld_vec_2;
    wire [23:0] in_chan_dep_data_vec_2;
    wire [1:0] token_in_vec_2;
    wire [1:0] out_chan_dep_vld_vec_2;
    wire [11:0] out_chan_dep_data_2;
    wire [1:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [11:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_6_2;
    wire [11:0] dep_chan_data_6_2;
    wire token_6_2;
    wire [1:0] proc_dep_vld_vec_3;
    reg [1:0] proc_dep_vld_vec_3_reg;
    wire [1:0] in_chan_dep_vld_vec_3;
    wire [23:0] in_chan_dep_data_vec_3;
    wire [1:0] token_in_vec_3;
    wire [1:0] out_chan_dep_vld_vec_3;
    wire [11:0] out_chan_dep_data_3;
    wire [1:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_0_3;
    wire [11:0] dep_chan_data_0_3;
    wire token_0_3;
    wire dep_chan_vld_5_3;
    wire [11:0] dep_chan_data_5_3;
    wire token_5_3;
    wire [1:0] proc_dep_vld_vec_4;
    reg [1:0] proc_dep_vld_vec_4_reg;
    wire [1:0] in_chan_dep_vld_vec_4;
    wire [23:0] in_chan_dep_data_vec_4;
    wire [1:0] token_in_vec_4;
    wire [1:0] out_chan_dep_vld_vec_4;
    wire [11:0] out_chan_dep_data_4;
    wire [1:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_0_4;
    wire [11:0] dep_chan_data_0_4;
    wire token_0_4;
    wire dep_chan_vld_6_4;
    wire [11:0] dep_chan_data_6_4;
    wire token_6_4;
    wire [3:0] proc_dep_vld_vec_5;
    reg [3:0] proc_dep_vld_vec_5_reg;
    wire [3:0] in_chan_dep_vld_vec_5;
    wire [47:0] in_chan_dep_data_vec_5;
    wire [3:0] token_in_vec_5;
    wire [3:0] out_chan_dep_vld_vec_5;
    wire [11:0] out_chan_dep_data_5;
    wire [3:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_1_5;
    wire [11:0] dep_chan_data_1_5;
    wire token_1_5;
    wire dep_chan_vld_3_5;
    wire [11:0] dep_chan_data_3_5;
    wire token_3_5;
    wire dep_chan_vld_7_5;
    wire [11:0] dep_chan_data_7_5;
    wire token_7_5;
    wire dep_chan_vld_9_5;
    wire [11:0] dep_chan_data_9_5;
    wire token_9_5;
    wire [3:0] proc_dep_vld_vec_6;
    reg [3:0] proc_dep_vld_vec_6_reg;
    wire [3:0] in_chan_dep_vld_vec_6;
    wire [47:0] in_chan_dep_data_vec_6;
    wire [3:0] token_in_vec_6;
    wire [3:0] out_chan_dep_vld_vec_6;
    wire [11:0] out_chan_dep_data_6;
    wire [3:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_2_6;
    wire [11:0] dep_chan_data_2_6;
    wire token_2_6;
    wire dep_chan_vld_4_6;
    wire [11:0] dep_chan_data_4_6;
    wire token_4_6;
    wire dep_chan_vld_8_6;
    wire [11:0] dep_chan_data_8_6;
    wire token_8_6;
    wire dep_chan_vld_10_6;
    wire [11:0] dep_chan_data_10_6;
    wire token_10_6;
    wire [0:0] proc_dep_vld_vec_7;
    reg [0:0] proc_dep_vld_vec_7_reg;
    wire [1:0] in_chan_dep_vld_vec_7;
    wire [23:0] in_chan_dep_data_vec_7;
    wire [1:0] token_in_vec_7;
    wire [0:0] out_chan_dep_vld_vec_7;
    wire [11:0] out_chan_dep_data_7;
    wire [0:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_5_7;
    wire [11:0] dep_chan_data_5_7;
    wire token_5_7;
    wire dep_chan_vld_9_7;
    wire [11:0] dep_chan_data_9_7;
    wire token_9_7;
    wire [0:0] proc_dep_vld_vec_8;
    reg [0:0] proc_dep_vld_vec_8_reg;
    wire [1:0] in_chan_dep_vld_vec_8;
    wire [23:0] in_chan_dep_data_vec_8;
    wire [1:0] token_in_vec_8;
    wire [0:0] out_chan_dep_vld_vec_8;
    wire [11:0] out_chan_dep_data_8;
    wire [0:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_6_8;
    wire [11:0] dep_chan_data_6_8;
    wire token_6_8;
    wire dep_chan_vld_10_8;
    wire [11:0] dep_chan_data_10_8;
    wire token_10_8;
    wire [2:0] proc_dep_vld_vec_9;
    reg [2:0] proc_dep_vld_vec_9_reg;
    wire [1:0] in_chan_dep_vld_vec_9;
    wire [23:0] in_chan_dep_data_vec_9;
    wire [1:0] token_in_vec_9;
    wire [2:0] out_chan_dep_vld_vec_9;
    wire [11:0] out_chan_dep_data_9;
    wire [2:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_5_9;
    wire [11:0] dep_chan_data_5_9;
    wire token_5_9;
    wire dep_chan_vld_11_9;
    wire [11:0] dep_chan_data_11_9;
    wire token_11_9;
    wire [2:0] proc_dep_vld_vec_10;
    reg [2:0] proc_dep_vld_vec_10_reg;
    wire [1:0] in_chan_dep_vld_vec_10;
    wire [23:0] in_chan_dep_data_vec_10;
    wire [1:0] token_in_vec_10;
    wire [2:0] out_chan_dep_vld_vec_10;
    wire [11:0] out_chan_dep_data_10;
    wire [2:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_6_10;
    wire [11:0] dep_chan_data_6_10;
    wire token_6_10;
    wire dep_chan_vld_11_10;
    wire [11:0] dep_chan_data_11_10;
    wire token_11_10;
    wire [1:0] proc_dep_vld_vec_11;
    reg [1:0] proc_dep_vld_vec_11_reg;
    wire [1:0] in_chan_dep_vld_vec_11;
    wire [23:0] in_chan_dep_data_vec_11;
    wire [1:0] token_in_vec_11;
    wire [1:0] out_chan_dep_vld_vec_11;
    wire [11:0] out_chan_dep_data_11;
    wire [1:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_9_11;
    wire [11:0] dep_chan_data_9_11;
    wire token_9_11;
    wire dep_chan_vld_10_11;
    wire [11:0] dep_chan_data_10_11;
    wire token_10_11;
    wire [11:0] dl_in_vec;
    wire dl_detect_out;
    wire [11:0] origin;
    wire token_clear;

    reg ap_done_reg_0;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_done;
        end
    end

    reg ap_done_reg_1;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_done;
        end
    end

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0
    AESL_deadlock_detect_unit #(12, 0, 4, 4) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0.data_q_V_out_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.ap_done));
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0.data_q_V_out1_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.ap_done));
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0.data_vk_V_out_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.ap_done));
    assign proc_dep_vld_vec_0[3] = dl_detect_out ? proc_dep_vld_vec_0_reg[3] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.multiheadattention_ap_fixed_ap_fixed_33_13_5_3_0_config3_entry333_U0.data_vk_V_out2_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.ap_done));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[11 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[23 : 12] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_3_0;
    assign in_chan_dep_data_vec_0[35 : 24] = dep_chan_data_3_0;
    assign token_in_vec_0[2] = token_3_0;
    assign in_chan_dep_vld_vec_0[3] = dep_chan_vld_4_0;
    assign in_chan_dep_data_vec_0[47 : 36] = dep_chan_data_4_0;
    assign token_in_vec_0[3] = token_4_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[1];
    assign dep_chan_vld_0_3 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_3 = out_chan_dep_data_0;
    assign token_0_3 = token_out_vec_0[2];
    assign dep_chan_vld_0_4 = out_chan_dep_vld_vec_0[3];
    assign dep_chan_data_0_4 = out_chan_dep_data_0;
    assign token_0_4 = token_out_vec_0[3];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0
    AESL_deadlock_detect_unit #(12, 1, 2, 2) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.data_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0$ap_idle)));
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.d_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.d_V_V1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.d_V_V2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_166_U0.d_V_V3_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170hbi_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.ap_done));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[11 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_5_1;
    assign in_chan_dep_data_vec_1[23 : 12] = dep_chan_data_5_1;
    assign token_in_vec_1[1] = token_5_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];
    assign dep_chan_vld_1_5 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_5 = out_chan_dep_data_1;
    assign token_1_5 = token_out_vec_1[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0
    AESL_deadlock_detect_unit #(12, 2, 2, 2) AESL_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.data_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0$ap_idle)));
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.d_V_V14_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.d_V_V15_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.d_V_V16_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_167_U0.d_V_V17_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171ibs_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.ap_done));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[11 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_6_2;
    assign in_chan_dep_data_vec_2[23 : 12] = dep_chan_data_6_2;
    assign token_in_vec_2[1] = token_6_2;
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[0];
    assign dep_chan_vld_2_6 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_6 = out_chan_dep_data_2;
    assign token_2_6 = token_out_vec_2[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0
    AESL_deadlock_detect_unit #(12, 3, 2, 2) AESL_deadlock_detect_unit_3 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.data_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0$ap_idle)));
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.d_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.d_V_V1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.d_V_V2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_168_U0.d_V_V3_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_0_3;
    assign in_chan_dep_data_vec_3[11 : 0] = dep_chan_data_0_3;
    assign token_in_vec_3[0] = token_0_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_5_3;
    assign in_chan_dep_data_vec_3[23 : 12] = dep_chan_data_5_3;
    assign token_in_vec_3[1] = token_5_3;
    assign dep_chan_vld_3_0 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_0 = out_chan_dep_data_3;
    assign token_3_0 = token_out_vec_3[0];
    assign dep_chan_vld_3_5 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_5 = out_chan_dep_data_3;
    assign token_3_5 = token_out_vec_3[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0
    AESL_deadlock_detect_unit #(12, 4, 2, 2) AESL_deadlock_detect_unit_4 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.data_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0$ap_idle)));
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.d_V_V14_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.d_V_V15_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.d_V_V16_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.data_prep_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_169_U0.d_V_V17_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_0_4;
    assign in_chan_dep_data_vec_4[11 : 0] = dep_chan_data_0_4;
    assign token_in_vec_4[0] = token_0_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_6_4;
    assign in_chan_dep_data_vec_4[23 : 12] = dep_chan_data_6_4;
    assign token_in_vec_4[1] = token_6_4;
    assign dep_chan_vld_4_0 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_0 = out_chan_dep_data_4;
    assign token_4_0 = token_out_vec_4[0];
    assign dep_chan_vld_4_6 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_6 = out_chan_dep_data_4;
    assign token_4_6 = token_out_vec_4[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0
    AESL_deadlock_detect_unit #(12, 5, 4, 4) AESL_deadlock_detect_unit_5 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_0_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_1_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_2_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_3_V_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170hbi_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0$ap_idle)));
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_0_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_1_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_2_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_3_V_V_blk_n);
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.k_proj_V_data_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.q_proj_V_data_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0.ap_done));
    assign proc_dep_vld_vec_5[3] = dl_detect_out ? proc_dep_vld_vec_5_reg[3] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_170_U0.v_proj_V_data_V_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_1_5;
    assign in_chan_dep_data_vec_5[11 : 0] = dep_chan_data_1_5;
    assign token_in_vec_5[0] = token_1_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_3_5;
    assign in_chan_dep_data_vec_5[23 : 12] = dep_chan_data_3_5;
    assign token_in_vec_5[1] = token_3_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_7_5;
    assign in_chan_dep_data_vec_5[35 : 24] = dep_chan_data_7_5;
    assign token_in_vec_5[2] = token_7_5;
    assign in_chan_dep_vld_vec_5[3] = dep_chan_vld_9_5;
    assign in_chan_dep_data_vec_5[47 : 36] = dep_chan_data_9_5;
    assign token_in_vec_5[3] = token_9_5;
    assign dep_chan_vld_5_1 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_1 = out_chan_dep_data_5;
    assign token_5_1 = token_out_vec_5[0];
    assign dep_chan_vld_5_3 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_3 = out_chan_dep_data_5;
    assign token_5_3 = token_out_vec_5[1];
    assign dep_chan_vld_5_7 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_7 = out_chan_dep_data_5;
    assign token_5_7 = token_out_vec_5[2];
    assign dep_chan_vld_5_9 = out_chan_dep_vld_vec_5[3];
    assign dep_chan_data_5_9 = out_chan_dep_data_5;
    assign token_5_9 = token_out_vec_5[3];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0
    AESL_deadlock_detect_unit #(12, 6, 4, 4) AESL_deadlock_detect_unit_6 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_0_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_1_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_2_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_113.data_in_3_V_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171ibs_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0$ap_idle)));
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_0_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_1_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_2_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_125.data_in_3_V_V_blk_n);
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.k_proj_V_data_V3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.q_proj_V_data_V4_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0.ap_done));
    assign proc_dep_vld_vec_6[3] = dl_detect_out ? proc_dep_vld_vec_6_reg[3] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.lin_projection_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_171_U0.v_proj_V_data_V5_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_2_6;
    assign in_chan_dep_data_vec_6[11 : 0] = dep_chan_data_2_6;
    assign token_in_vec_6[0] = token_2_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_4_6;
    assign in_chan_dep_data_vec_6[23 : 12] = dep_chan_data_4_6;
    assign token_in_vec_6[1] = token_4_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_8_6;
    assign in_chan_dep_data_vec_6[35 : 24] = dep_chan_data_8_6;
    assign token_in_vec_6[2] = token_8_6;
    assign in_chan_dep_vld_vec_6[3] = dep_chan_vld_10_6;
    assign in_chan_dep_data_vec_6[47 : 36] = dep_chan_data_10_6;
    assign token_in_vec_6[3] = token_10_6;
    assign dep_chan_vld_6_2 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_2 = out_chan_dep_data_6;
    assign token_6_2 = token_out_vec_6[0];
    assign dep_chan_vld_6_4 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_4 = out_chan_dep_data_6;
    assign token_6_4 = token_out_vec_6[1];
    assign dep_chan_vld_6_8 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_8 = out_chan_dep_data_6;
    assign token_6_8 = token_out_vec_6[2];
    assign dep_chan_vld_6_10 = out_chan_dep_vld_vec_6[3];
    assign dep_chan_data_6_10 = out_chan_dep_data_6;
    assign token_6_10 = token_out_vec_6[3];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0
    AESL_deadlock_detect_unit #(12, 7, 2, 1) AESL_deadlock_detect_unit_7 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0.Q_V_data_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0.K_V_data_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_172_U0$ap_idle)));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_5_7;
    assign in_chan_dep_data_vec_7[11 : 0] = dep_chan_data_5_7;
    assign token_in_vec_7[0] = token_5_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_9_7;
    assign in_chan_dep_data_vec_7[23 : 12] = dep_chan_data_9_7;
    assign token_in_vec_7[1] = token_9_7;
    assign dep_chan_vld_7_5 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_5 = out_chan_dep_data_7;
    assign token_7_5 = token_out_vec_7[0];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0
    AESL_deadlock_detect_unit #(12, 8, 2, 1) AESL_deadlock_detect_unit_8 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0.Q_V_data_V1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0.K_V_data_V2_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_transpose_ap_fixed_ap_fixed_33_13_5_3_0_config3_173_U0$ap_idle)));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_6_8;
    assign in_chan_dep_data_vec_8[11 : 0] = dep_chan_data_6_8;
    assign token_in_vec_8[0] = token_6_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_10_8;
    assign in_chan_dep_data_vec_8[23 : 12] = dep_chan_data_10_8;
    assign token_in_vec_8[1] = token_10_8;
    assign dep_chan_vld_8_6 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_6 = out_chan_dep_data_8;
    assign token_8_6 = token_out_vec_8[0];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0
    AESL_deadlock_detect_unit #(12, 9, 2, 3) AESL_deadlock_detect_unit_9 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_0_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_1_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_2_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_3_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_4_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_5_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_6_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_7_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_8_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_9_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_10_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_11_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_12_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_13_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_14_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_15_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_16_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_17_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_18_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_0_19_19_V_U.if_write);
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.V_V_data_V_blk_n);
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.S_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_174_U0.S_V_V40_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_full_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_done));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_5_9;
    assign in_chan_dep_data_vec_9[11 : 0] = dep_chan_data_5_9;
    assign token_in_vec_9[0] = token_5_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_11_9;
    assign in_chan_dep_data_vec_9[23 : 12] = dep_chan_data_11_9;
    assign token_in_vec_9[1] = token_11_9;
    assign dep_chan_vld_9_7 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_7 = out_chan_dep_data_9;
    assign token_9_7 = token_out_vec_9[0];
    assign dep_chan_vld_9_5 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_5 = out_chan_dep_data_9;
    assign token_9_5 = token_out_vec_9[1];
    assign dep_chan_vld_9_11 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_11 = out_chan_dep_data_9;
    assign token_9_11 = token_out_vec_9[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0
    AESL_deadlock_detect_unit #(12, 10, 2, 3) AESL_deadlock_detect_unit_10 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_0_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_1_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_2_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_3_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_4_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_5_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_6_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_7_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_8_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_9_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_10_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_11_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_12_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_13_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_14_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_15_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_16_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_17_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_18_19_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_0_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_0_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_1_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_1_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_2_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_2_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_3_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_3_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_4_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_4_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_5_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_5_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_6_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_6_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_7_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_7_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_8_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_8_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_9_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_9_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_10_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_10_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_11_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_11_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_12_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_12_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_13_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_13_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_14_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_14_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_15_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_15_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_16_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_16_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_17_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_17_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_18_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_18_V_U.if_write | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_19_V_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_ready | AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.ap_idle) & ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.qk_mul_1_19_19_V_U.if_write);
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.V_V_data_V2_blk_n);
    assign proc_dep_vld_vec_10[2] = dl_detect_out ? proc_dep_vld_vec_10_reg[2] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.S_V_V3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.matrixmul_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_175_U0.S_V_V341_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_6_10;
    assign in_chan_dep_data_vec_10[11 : 0] = dep_chan_data_6_10;
    assign token_in_vec_10[0] = token_6_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_11_10;
    assign in_chan_dep_data_vec_10[23 : 12] = dep_chan_data_11_10;
    assign token_in_vec_10[1] = token_11_10;
    assign dep_chan_vld_10_8 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_8 = out_chan_dep_data_10;
    assign token_10_8 = token_out_vec_10[0];
    assign dep_chan_vld_10_6 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_6 = out_chan_dep_data_10;
    assign token_10_6 = token_out_vec_10[1];
    assign dep_chan_vld_10_11 = out_chan_dep_vld_vec_10[2];
    assign dep_chan_data_10_11 = out_chan_dep_data_10;
    assign token_10_11 = token_out_vec_10[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0$ap_idle <= AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0
    AESL_deadlock_detect_unit #(12, 11, 2, 2) AESL_deadlock_detect_unit_11 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.data_in_0_0_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.data_in_0_1_V_V_blk_n | (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.start_for_dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0_U.if_empty_n & (AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.ap_ready | AESL_inst_myproject$grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196$dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0$ap_idle)));
    assign proc_dep_vld_vec_11[1] = dl_detect_out ? proc_dep_vld_vec_11_reg[1] : (~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.data_in_1_0_V_V_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_16_6_5_3_0_ap_fixed_33_13_5_3_0_config3_s_fu_196.dense_out_ap_fixed_33_13_5_3_0_ap_fixed_33_13_5_3_0_config3_U0.data_in_1_1_V_V_blk_n);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_9_11;
    assign in_chan_dep_data_vec_11[11 : 0] = dep_chan_data_9_11;
    assign token_in_vec_11[0] = token_9_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_10_11;
    assign in_chan_dep_data_vec_11[23 : 12] = dep_chan_data_10_11;
    assign token_in_vec_11[1] = token_10_11;
    assign dep_chan_vld_11_9 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_9 = out_chan_dep_data_11;
    assign token_11_9 = token_out_vec_11[0];
    assign dep_chan_vld_11_10 = out_chan_dep_vld_vec_11[1];
    assign dep_chan_data_11_10 = out_chan_dep_data_11;
    assign token_11_10 = token_out_vec_11[1];


    AESL_deadlock_report_unit #(12) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
