
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_0_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_0_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_0_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_1_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_1_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_1_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_1_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_1_blk_n);
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_2_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_2_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_2_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_2_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_2_blk_n);
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_3_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_3_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_3_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_3_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_3_blk_n);
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_4_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_4_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_0_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_0_blk_n);
    assign fifo_intf_5.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_0_blk_n);
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_5_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_5_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_1_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_1_blk_n);
    assign fifo_intf_6.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_1_blk_n);
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_6_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_6_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_2_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_2_blk_n);
    assign fifo_intf_7.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_2_blk_n);
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_7_U.if_empty_n;
    assign fifo_intf_8.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_query_7_U.if_full_n;
    assign fifo_intf_8.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_3_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_3_blk_n);
    assign fifo_intf_8.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_3_blk_n);
    assign fifo_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_U.if_empty_n;
    assign fifo_intf_9.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_U.if_full_n;
    assign fifo_intf_9.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_0_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_0_blk_n);
    assign fifo_intf_9.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_0_blk_n);
    assign fifo_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_1_U.if_empty_n;
    assign fifo_intf_10.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_1_U.if_full_n;
    assign fifo_intf_10.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_1_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_1_blk_n);
    assign fifo_intf_10.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_1_blk_n);
    assign fifo_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_2_U.if_empty_n;
    assign fifo_intf_11.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_2_U.if_full_n;
    assign fifo_intf_11.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_2_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_2_blk_n);
    assign fifo_intf_11.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_2_blk_n);
    assign fifo_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_3_U.if_empty_n;
    assign fifo_intf_12.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_3_U.if_full_n;
    assign fifo_intf_12.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_3_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_3_blk_n);
    assign fifo_intf_12.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_3_blk_n);
    assign fifo_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_4_U.if_empty_n;
    assign fifo_intf_13.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_4_U.if_full_n;
    assign fifo_intf_13.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_0_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_0_blk_n);
    assign fifo_intf_13.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_0_blk_n);
    assign fifo_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_5_U.if_empty_n;
    assign fifo_intf_14.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_5_U.if_full_n;
    assign fifo_intf_14.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_1_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_1_blk_n);
    assign fifo_intf_14.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_1_blk_n);
    assign fifo_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_6_U.if_empty_n;
    assign fifo_intf_15.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_6_U.if_full_n;
    assign fifo_intf_15.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_2_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_2_blk_n);
    assign fifo_intf_15.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_2_blk_n);
    assign fifo_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_7_U.if_empty_n;
    assign fifo_intf_16.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.d_value_7_U.if_full_n;
    assign fifo_intf_16.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_3_blk_n & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_3_blk_n);
    assign fifo_intf_16.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_3_blk_n);
    assign fifo_intf_16.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_0_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_0_U.if_empty_n;
    assign fifo_intf_17.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_0_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_0_U.if_full_n;
    assign fifo_intf_17.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.k_proj_0_blk_n);
    assign fifo_intf_17.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.k_proj_0_blk_n);
    assign fifo_intf_17.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_0_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_0_U.if_empty_n;
    assign fifo_intf_18.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_0_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_0_U.if_full_n;
    assign fifo_intf_18.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.q_proj_0_blk_n);
    assign fifo_intf_18.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.q_proj_0_blk_n);
    assign fifo_intf_18.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_0_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_0_U.if_empty_n;
    assign fifo_intf_19.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_0_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_0_U.if_full_n;
    assign fifo_intf_19.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.v_proj_0_blk_n);
    assign fifo_intf_19.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.v_proj_0_blk_n);
    assign fifo_intf_19.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_1_U.if_empty_n;
    assign fifo_intf_20.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.k_proj_1_U.if_full_n;
    assign fifo_intf_20.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.k_proj_1_blk_n);
    assign fifo_intf_20.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.k_proj_1_blk_n);
    assign fifo_intf_20.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_1_U.if_empty_n;
    assign fifo_intf_21.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.q_proj_1_U.if_full_n;
    assign fifo_intf_21.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.q_proj_1_blk_n);
    assign fifo_intf_21.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.q_proj_1_blk_n);
    assign fifo_intf_21.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_1_U.if_empty_n;
    assign fifo_intf_22.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.v_proj_1_U.if_full_n;
    assign fifo_intf_22.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.v_proj_1_blk_n);
    assign fifo_intf_22.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.v_proj_1_blk_n);
    assign fifo_intf_22.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_U.if_empty_n;
    assign fifo_intf_23.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_U.if_full_n;
    assign fifo_intf_23.fifo_rd_block = 0;
    assign fifo_intf_23.fifo_wr_block = 0;
    assign fifo_intf_23.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_U.if_empty_n;
    assign fifo_intf_24.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_U.if_full_n;
    assign fifo_intf_24.fifo_rd_block = 0;
    assign fifo_intf_24.fifo_wr_block = 0;
    assign fifo_intf_24.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_U.if_empty_n;
    assign fifo_intf_25.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_U.if_full_n;
    assign fifo_intf_25.fifo_rd_block = 0;
    assign fifo_intf_25.fifo_wr_block = 0;
    assign fifo_intf_25.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_U.if_empty_n;
    assign fifo_intf_26.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_U.if_full_n;
    assign fifo_intf_26.fifo_rd_block = 0;
    assign fifo_intf_26.fifo_wr_block = 0;
    assign fifo_intf_26.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_U.if_empty_n;
    assign fifo_intf_27.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_U.if_full_n;
    assign fifo_intf_27.fifo_rd_block = 0;
    assign fifo_intf_27.fifo_wr_block = 0;
    assign fifo_intf_27.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_U.if_empty_n;
    assign fifo_intf_28.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_U.if_full_n;
    assign fifo_intf_28.fifo_rd_block = 0;
    assign fifo_intf_28.fifo_wr_block = 0;
    assign fifo_intf_28.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_U.if_empty_n;
    assign fifo_intf_29.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_U.if_full_n;
    assign fifo_intf_29.fifo_rd_block = 0;
    assign fifo_intf_29.fifo_wr_block = 0;
    assign fifo_intf_29.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_U.if_empty_n;
    assign fifo_intf_30.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_U.if_full_n;
    assign fifo_intf_30.fifo_rd_block = 0;
    assign fifo_intf_30.fifo_wr_block = 0;
    assign fifo_intf_30.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_U.if_empty_n;
    assign fifo_intf_31.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_U.if_full_n;
    assign fifo_intf_31.fifo_rd_block = 0;
    assign fifo_intf_31.fifo_wr_block = 0;
    assign fifo_intf_31.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_U.if_empty_n;
    assign fifo_intf_32.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_U.if_full_n;
    assign fifo_intf_32.fifo_rd_block = 0;
    assign fifo_intf_32.fifo_wr_block = 0;
    assign fifo_intf_32.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_U.if_empty_n;
    assign fifo_intf_33.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_U.if_full_n;
    assign fifo_intf_33.fifo_rd_block = 0;
    assign fifo_intf_33.fifo_wr_block = 0;
    assign fifo_intf_33.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_U.if_empty_n;
    assign fifo_intf_34.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_U.if_full_n;
    assign fifo_intf_34.fifo_rd_block = 0;
    assign fifo_intf_34.fifo_wr_block = 0;
    assign fifo_intf_34.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;
    df_fifo_intf fifo_intf_35(clock,reset);
    assign fifo_intf_35.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_U.if_empty_n;
    assign fifo_intf_35.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_U.if_full_n;
    assign fifo_intf_35.fifo_rd_block = 0;
    assign fifo_intf_35.fifo_wr_block = 0;
    assign fifo_intf_35.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_35;
    csv_file_dump cstatus_csv_dumper_35;
    df_fifo_monitor fifo_monitor_35;
    df_fifo_intf fifo_intf_36(clock,reset);
    assign fifo_intf_36.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_U.if_empty_n;
    assign fifo_intf_36.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_U.if_full_n;
    assign fifo_intf_36.fifo_rd_block = 0;
    assign fifo_intf_36.fifo_wr_block = 0;
    assign fifo_intf_36.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_36;
    csv_file_dump cstatus_csv_dumper_36;
    df_fifo_monitor fifo_monitor_36;
    df_fifo_intf fifo_intf_37(clock,reset);
    assign fifo_intf_37.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_U.if_empty_n;
    assign fifo_intf_37.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_U.if_full_n;
    assign fifo_intf_37.fifo_rd_block = 0;
    assign fifo_intf_37.fifo_wr_block = 0;
    assign fifo_intf_37.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_37;
    csv_file_dump cstatus_csv_dumper_37;
    df_fifo_monitor fifo_monitor_37;
    df_fifo_intf fifo_intf_38(clock,reset);
    assign fifo_intf_38.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_U.if_empty_n;
    assign fifo_intf_38.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_U.if_full_n;
    assign fifo_intf_38.fifo_rd_block = 0;
    assign fifo_intf_38.fifo_wr_block = 0;
    assign fifo_intf_38.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_38;
    csv_file_dump cstatus_csv_dumper_38;
    df_fifo_monitor fifo_monitor_38;
    df_fifo_intf fifo_intf_39(clock,reset);
    assign fifo_intf_39.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_U.if_empty_n;
    assign fifo_intf_39.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_U.if_full_n;
    assign fifo_intf_39.fifo_rd_block = 0;
    assign fifo_intf_39.fifo_wr_block = 0;
    assign fifo_intf_39.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_39;
    csv_file_dump cstatus_csv_dumper_39;
    df_fifo_monitor fifo_monitor_39;
    df_fifo_intf fifo_intf_40(clock,reset);
    assign fifo_intf_40.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_U.if_empty_n;
    assign fifo_intf_40.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_U.if_full_n;
    assign fifo_intf_40.fifo_rd_block = 0;
    assign fifo_intf_40.fifo_wr_block = 0;
    assign fifo_intf_40.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_40;
    csv_file_dump cstatus_csv_dumper_40;
    df_fifo_monitor fifo_monitor_40;
    df_fifo_intf fifo_intf_41(clock,reset);
    assign fifo_intf_41.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_U.if_empty_n;
    assign fifo_intf_41.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_U.if_full_n;
    assign fifo_intf_41.fifo_rd_block = 0;
    assign fifo_intf_41.fifo_wr_block = 0;
    assign fifo_intf_41.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_41;
    csv_file_dump cstatus_csv_dumper_41;
    df_fifo_monitor fifo_monitor_41;
    df_fifo_intf fifo_intf_42(clock,reset);
    assign fifo_intf_42.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_U.if_empty_n;
    assign fifo_intf_42.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_U.if_full_n;
    assign fifo_intf_42.fifo_rd_block = 0;
    assign fifo_intf_42.fifo_wr_block = 0;
    assign fifo_intf_42.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_42;
    csv_file_dump cstatus_csv_dumper_42;
    df_fifo_monitor fifo_monitor_42;
    df_fifo_intf fifo_intf_43(clock,reset);
    assign fifo_intf_43.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_1_U.if_empty_n;
    assign fifo_intf_43.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_1_U.if_full_n;
    assign fifo_intf_43.fifo_rd_block = 0;
    assign fifo_intf_43.fifo_wr_block = 0;
    assign fifo_intf_43.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_43;
    csv_file_dump cstatus_csv_dumper_43;
    df_fifo_monitor fifo_monitor_43;
    df_fifo_intf fifo_intf_44(clock,reset);
    assign fifo_intf_44.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_1_U.if_empty_n;
    assign fifo_intf_44.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_1_U.if_full_n;
    assign fifo_intf_44.fifo_rd_block = 0;
    assign fifo_intf_44.fifo_wr_block = 0;
    assign fifo_intf_44.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_44;
    csv_file_dump cstatus_csv_dumper_44;
    df_fifo_monitor fifo_monitor_44;
    df_fifo_intf fifo_intf_45(clock,reset);
    assign fifo_intf_45.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_1_U.if_empty_n;
    assign fifo_intf_45.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_1_U.if_full_n;
    assign fifo_intf_45.fifo_rd_block = 0;
    assign fifo_intf_45.fifo_wr_block = 0;
    assign fifo_intf_45.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_45;
    csv_file_dump cstatus_csv_dumper_45;
    df_fifo_monitor fifo_monitor_45;
    df_fifo_intf fifo_intf_46(clock,reset);
    assign fifo_intf_46.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_1_U.if_empty_n;
    assign fifo_intf_46.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_1_U.if_full_n;
    assign fifo_intf_46.fifo_rd_block = 0;
    assign fifo_intf_46.fifo_wr_block = 0;
    assign fifo_intf_46.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_46;
    csv_file_dump cstatus_csv_dumper_46;
    df_fifo_monitor fifo_monitor_46;
    df_fifo_intf fifo_intf_47(clock,reset);
    assign fifo_intf_47.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_1_U.if_empty_n;
    assign fifo_intf_47.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_1_U.if_full_n;
    assign fifo_intf_47.fifo_rd_block = 0;
    assign fifo_intf_47.fifo_wr_block = 0;
    assign fifo_intf_47.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_47;
    csv_file_dump cstatus_csv_dumper_47;
    df_fifo_monitor fifo_monitor_47;
    df_fifo_intf fifo_intf_48(clock,reset);
    assign fifo_intf_48.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_1_U.if_empty_n;
    assign fifo_intf_48.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_1_U.if_full_n;
    assign fifo_intf_48.fifo_rd_block = 0;
    assign fifo_intf_48.fifo_wr_block = 0;
    assign fifo_intf_48.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_48;
    csv_file_dump cstatus_csv_dumper_48;
    df_fifo_monitor fifo_monitor_48;
    df_fifo_intf fifo_intf_49(clock,reset);
    assign fifo_intf_49.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_1_U.if_empty_n;
    assign fifo_intf_49.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_1_U.if_full_n;
    assign fifo_intf_49.fifo_rd_block = 0;
    assign fifo_intf_49.fifo_wr_block = 0;
    assign fifo_intf_49.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_49;
    csv_file_dump cstatus_csv_dumper_49;
    df_fifo_monitor fifo_monitor_49;
    df_fifo_intf fifo_intf_50(clock,reset);
    assign fifo_intf_50.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_1_U.if_empty_n;
    assign fifo_intf_50.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_1_U.if_full_n;
    assign fifo_intf_50.fifo_rd_block = 0;
    assign fifo_intf_50.fifo_wr_block = 0;
    assign fifo_intf_50.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_50;
    csv_file_dump cstatus_csv_dumper_50;
    df_fifo_monitor fifo_monitor_50;
    df_fifo_intf fifo_intf_51(clock,reset);
    assign fifo_intf_51.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_1_U.if_empty_n;
    assign fifo_intf_51.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_1_U.if_full_n;
    assign fifo_intf_51.fifo_rd_block = 0;
    assign fifo_intf_51.fifo_wr_block = 0;
    assign fifo_intf_51.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_51;
    csv_file_dump cstatus_csv_dumper_51;
    df_fifo_monitor fifo_monitor_51;
    df_fifo_intf fifo_intf_52(clock,reset);
    assign fifo_intf_52.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_1_U.if_empty_n;
    assign fifo_intf_52.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_1_U.if_full_n;
    assign fifo_intf_52.fifo_rd_block = 0;
    assign fifo_intf_52.fifo_wr_block = 0;
    assign fifo_intf_52.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_52;
    csv_file_dump cstatus_csv_dumper_52;
    df_fifo_monitor fifo_monitor_52;
    df_fifo_intf fifo_intf_53(clock,reset);
    assign fifo_intf_53.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_1_U.if_empty_n;
    assign fifo_intf_53.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_1_U.if_full_n;
    assign fifo_intf_53.fifo_rd_block = 0;
    assign fifo_intf_53.fifo_wr_block = 0;
    assign fifo_intf_53.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_53;
    csv_file_dump cstatus_csv_dumper_53;
    df_fifo_monitor fifo_monitor_53;
    df_fifo_intf fifo_intf_54(clock,reset);
    assign fifo_intf_54.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_1_U.if_empty_n;
    assign fifo_intf_54.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_1_U.if_full_n;
    assign fifo_intf_54.fifo_rd_block = 0;
    assign fifo_intf_54.fifo_wr_block = 0;
    assign fifo_intf_54.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_54;
    csv_file_dump cstatus_csv_dumper_54;
    df_fifo_monitor fifo_monitor_54;
    df_fifo_intf fifo_intf_55(clock,reset);
    assign fifo_intf_55.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_1_U.if_empty_n;
    assign fifo_intf_55.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_1_U.if_full_n;
    assign fifo_intf_55.fifo_rd_block = 0;
    assign fifo_intf_55.fifo_wr_block = 0;
    assign fifo_intf_55.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_55;
    csv_file_dump cstatus_csv_dumper_55;
    df_fifo_monitor fifo_monitor_55;
    df_fifo_intf fifo_intf_56(clock,reset);
    assign fifo_intf_56.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_1_U.if_empty_n;
    assign fifo_intf_56.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_1_U.if_full_n;
    assign fifo_intf_56.fifo_rd_block = 0;
    assign fifo_intf_56.fifo_wr_block = 0;
    assign fifo_intf_56.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_56;
    csv_file_dump cstatus_csv_dumper_56;
    df_fifo_monitor fifo_monitor_56;
    df_fifo_intf fifo_intf_57(clock,reset);
    assign fifo_intf_57.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_1_U.if_empty_n;
    assign fifo_intf_57.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_1_U.if_full_n;
    assign fifo_intf_57.fifo_rd_block = 0;
    assign fifo_intf_57.fifo_wr_block = 0;
    assign fifo_intf_57.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_57;
    csv_file_dump cstatus_csv_dumper_57;
    df_fifo_monitor fifo_monitor_57;
    df_fifo_intf fifo_intf_58(clock,reset);
    assign fifo_intf_58.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_1_U.if_empty_n;
    assign fifo_intf_58.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_1_U.if_full_n;
    assign fifo_intf_58.fifo_rd_block = 0;
    assign fifo_intf_58.fifo_wr_block = 0;
    assign fifo_intf_58.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_58;
    csv_file_dump cstatus_csv_dumper_58;
    df_fifo_monitor fifo_monitor_58;
    df_fifo_intf fifo_intf_59(clock,reset);
    assign fifo_intf_59.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_1_U.if_empty_n;
    assign fifo_intf_59.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_1_U.if_full_n;
    assign fifo_intf_59.fifo_rd_block = 0;
    assign fifo_intf_59.fifo_wr_block = 0;
    assign fifo_intf_59.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_59;
    csv_file_dump cstatus_csv_dumper_59;
    df_fifo_monitor fifo_monitor_59;
    df_fifo_intf fifo_intf_60(clock,reset);
    assign fifo_intf_60.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_1_U.if_empty_n;
    assign fifo_intf_60.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_1_U.if_full_n;
    assign fifo_intf_60.fifo_rd_block = 0;
    assign fifo_intf_60.fifo_wr_block = 0;
    assign fifo_intf_60.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_60;
    csv_file_dump cstatus_csv_dumper_60;
    df_fifo_monitor fifo_monitor_60;
    df_fifo_intf fifo_intf_61(clock,reset);
    assign fifo_intf_61.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_1_U.if_empty_n;
    assign fifo_intf_61.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_1_U.if_full_n;
    assign fifo_intf_61.fifo_rd_block = 0;
    assign fifo_intf_61.fifo_wr_block = 0;
    assign fifo_intf_61.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_61;
    csv_file_dump cstatus_csv_dumper_61;
    df_fifo_monitor fifo_monitor_61;
    df_fifo_intf fifo_intf_62(clock,reset);
    assign fifo_intf_62.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_1_U.if_empty_n;
    assign fifo_intf_62.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_1_U.if_full_n;
    assign fifo_intf_62.fifo_rd_block = 0;
    assign fifo_intf_62.fifo_wr_block = 0;
    assign fifo_intf_62.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_62;
    csv_file_dump cstatus_csv_dumper_62;
    df_fifo_monitor fifo_monitor_62;
    df_fifo_intf fifo_intf_63(clock,reset);
    assign fifo_intf_63.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_2_U.if_empty_n;
    assign fifo_intf_63.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_2_U.if_full_n;
    assign fifo_intf_63.fifo_rd_block = 0;
    assign fifo_intf_63.fifo_wr_block = 0;
    assign fifo_intf_63.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_63;
    csv_file_dump cstatus_csv_dumper_63;
    df_fifo_monitor fifo_monitor_63;
    df_fifo_intf fifo_intf_64(clock,reset);
    assign fifo_intf_64.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_2_U.if_empty_n;
    assign fifo_intf_64.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_2_U.if_full_n;
    assign fifo_intf_64.fifo_rd_block = 0;
    assign fifo_intf_64.fifo_wr_block = 0;
    assign fifo_intf_64.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_64;
    csv_file_dump cstatus_csv_dumper_64;
    df_fifo_monitor fifo_monitor_64;
    df_fifo_intf fifo_intf_65(clock,reset);
    assign fifo_intf_65.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_2_U.if_empty_n;
    assign fifo_intf_65.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_2_U.if_full_n;
    assign fifo_intf_65.fifo_rd_block = 0;
    assign fifo_intf_65.fifo_wr_block = 0;
    assign fifo_intf_65.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_65;
    csv_file_dump cstatus_csv_dumper_65;
    df_fifo_monitor fifo_monitor_65;
    df_fifo_intf fifo_intf_66(clock,reset);
    assign fifo_intf_66.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_2_U.if_empty_n;
    assign fifo_intf_66.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_2_U.if_full_n;
    assign fifo_intf_66.fifo_rd_block = 0;
    assign fifo_intf_66.fifo_wr_block = 0;
    assign fifo_intf_66.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_66;
    csv_file_dump cstatus_csv_dumper_66;
    df_fifo_monitor fifo_monitor_66;
    df_fifo_intf fifo_intf_67(clock,reset);
    assign fifo_intf_67.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_2_U.if_empty_n;
    assign fifo_intf_67.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_2_U.if_full_n;
    assign fifo_intf_67.fifo_rd_block = 0;
    assign fifo_intf_67.fifo_wr_block = 0;
    assign fifo_intf_67.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_67;
    csv_file_dump cstatus_csv_dumper_67;
    df_fifo_monitor fifo_monitor_67;
    df_fifo_intf fifo_intf_68(clock,reset);
    assign fifo_intf_68.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_2_U.if_empty_n;
    assign fifo_intf_68.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_2_U.if_full_n;
    assign fifo_intf_68.fifo_rd_block = 0;
    assign fifo_intf_68.fifo_wr_block = 0;
    assign fifo_intf_68.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_68;
    csv_file_dump cstatus_csv_dumper_68;
    df_fifo_monitor fifo_monitor_68;
    df_fifo_intf fifo_intf_69(clock,reset);
    assign fifo_intf_69.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_2_U.if_empty_n;
    assign fifo_intf_69.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_2_U.if_full_n;
    assign fifo_intf_69.fifo_rd_block = 0;
    assign fifo_intf_69.fifo_wr_block = 0;
    assign fifo_intf_69.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_69;
    csv_file_dump cstatus_csv_dumper_69;
    df_fifo_monitor fifo_monitor_69;
    df_fifo_intf fifo_intf_70(clock,reset);
    assign fifo_intf_70.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_2_U.if_empty_n;
    assign fifo_intf_70.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_2_U.if_full_n;
    assign fifo_intf_70.fifo_rd_block = 0;
    assign fifo_intf_70.fifo_wr_block = 0;
    assign fifo_intf_70.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_70;
    csv_file_dump cstatus_csv_dumper_70;
    df_fifo_monitor fifo_monitor_70;
    df_fifo_intf fifo_intf_71(clock,reset);
    assign fifo_intf_71.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_2_U.if_empty_n;
    assign fifo_intf_71.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_2_U.if_full_n;
    assign fifo_intf_71.fifo_rd_block = 0;
    assign fifo_intf_71.fifo_wr_block = 0;
    assign fifo_intf_71.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_71;
    csv_file_dump cstatus_csv_dumper_71;
    df_fifo_monitor fifo_monitor_71;
    df_fifo_intf fifo_intf_72(clock,reset);
    assign fifo_intf_72.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_2_U.if_empty_n;
    assign fifo_intf_72.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_2_U.if_full_n;
    assign fifo_intf_72.fifo_rd_block = 0;
    assign fifo_intf_72.fifo_wr_block = 0;
    assign fifo_intf_72.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_72;
    csv_file_dump cstatus_csv_dumper_72;
    df_fifo_monitor fifo_monitor_72;
    df_fifo_intf fifo_intf_73(clock,reset);
    assign fifo_intf_73.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_2_U.if_empty_n;
    assign fifo_intf_73.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_2_U.if_full_n;
    assign fifo_intf_73.fifo_rd_block = 0;
    assign fifo_intf_73.fifo_wr_block = 0;
    assign fifo_intf_73.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_73;
    csv_file_dump cstatus_csv_dumper_73;
    df_fifo_monitor fifo_monitor_73;
    df_fifo_intf fifo_intf_74(clock,reset);
    assign fifo_intf_74.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_2_U.if_empty_n;
    assign fifo_intf_74.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_2_U.if_full_n;
    assign fifo_intf_74.fifo_rd_block = 0;
    assign fifo_intf_74.fifo_wr_block = 0;
    assign fifo_intf_74.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_74;
    csv_file_dump cstatus_csv_dumper_74;
    df_fifo_monitor fifo_monitor_74;
    df_fifo_intf fifo_intf_75(clock,reset);
    assign fifo_intf_75.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_2_U.if_empty_n;
    assign fifo_intf_75.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_2_U.if_full_n;
    assign fifo_intf_75.fifo_rd_block = 0;
    assign fifo_intf_75.fifo_wr_block = 0;
    assign fifo_intf_75.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_75;
    csv_file_dump cstatus_csv_dumper_75;
    df_fifo_monitor fifo_monitor_75;
    df_fifo_intf fifo_intf_76(clock,reset);
    assign fifo_intf_76.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_2_U.if_empty_n;
    assign fifo_intf_76.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_2_U.if_full_n;
    assign fifo_intf_76.fifo_rd_block = 0;
    assign fifo_intf_76.fifo_wr_block = 0;
    assign fifo_intf_76.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_76;
    csv_file_dump cstatus_csv_dumper_76;
    df_fifo_monitor fifo_monitor_76;
    df_fifo_intf fifo_intf_77(clock,reset);
    assign fifo_intf_77.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_2_U.if_empty_n;
    assign fifo_intf_77.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_2_U.if_full_n;
    assign fifo_intf_77.fifo_rd_block = 0;
    assign fifo_intf_77.fifo_wr_block = 0;
    assign fifo_intf_77.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_77;
    csv_file_dump cstatus_csv_dumper_77;
    df_fifo_monitor fifo_monitor_77;
    df_fifo_intf fifo_intf_78(clock,reset);
    assign fifo_intf_78.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_2_U.if_empty_n;
    assign fifo_intf_78.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_2_U.if_full_n;
    assign fifo_intf_78.fifo_rd_block = 0;
    assign fifo_intf_78.fifo_wr_block = 0;
    assign fifo_intf_78.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_78;
    csv_file_dump cstatus_csv_dumper_78;
    df_fifo_monitor fifo_monitor_78;
    df_fifo_intf fifo_intf_79(clock,reset);
    assign fifo_intf_79.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_2_U.if_empty_n;
    assign fifo_intf_79.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_2_U.if_full_n;
    assign fifo_intf_79.fifo_rd_block = 0;
    assign fifo_intf_79.fifo_wr_block = 0;
    assign fifo_intf_79.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_79;
    csv_file_dump cstatus_csv_dumper_79;
    df_fifo_monitor fifo_monitor_79;
    df_fifo_intf fifo_intf_80(clock,reset);
    assign fifo_intf_80.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_2_U.if_empty_n;
    assign fifo_intf_80.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_2_U.if_full_n;
    assign fifo_intf_80.fifo_rd_block = 0;
    assign fifo_intf_80.fifo_wr_block = 0;
    assign fifo_intf_80.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_80;
    csv_file_dump cstatus_csv_dumper_80;
    df_fifo_monitor fifo_monitor_80;
    df_fifo_intf fifo_intf_81(clock,reset);
    assign fifo_intf_81.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_2_U.if_empty_n;
    assign fifo_intf_81.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_2_U.if_full_n;
    assign fifo_intf_81.fifo_rd_block = 0;
    assign fifo_intf_81.fifo_wr_block = 0;
    assign fifo_intf_81.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_81;
    csv_file_dump cstatus_csv_dumper_81;
    df_fifo_monitor fifo_monitor_81;
    df_fifo_intf fifo_intf_82(clock,reset);
    assign fifo_intf_82.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_2_U.if_empty_n;
    assign fifo_intf_82.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_2_U.if_full_n;
    assign fifo_intf_82.fifo_rd_block = 0;
    assign fifo_intf_82.fifo_wr_block = 0;
    assign fifo_intf_82.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_82;
    csv_file_dump cstatus_csv_dumper_82;
    df_fifo_monitor fifo_monitor_82;
    df_fifo_intf fifo_intf_83(clock,reset);
    assign fifo_intf_83.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_3_U.if_empty_n;
    assign fifo_intf_83.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_3_U.if_full_n;
    assign fifo_intf_83.fifo_rd_block = 0;
    assign fifo_intf_83.fifo_wr_block = 0;
    assign fifo_intf_83.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_83;
    csv_file_dump cstatus_csv_dumper_83;
    df_fifo_monitor fifo_monitor_83;
    df_fifo_intf fifo_intf_84(clock,reset);
    assign fifo_intf_84.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_3_U.if_empty_n;
    assign fifo_intf_84.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_3_U.if_full_n;
    assign fifo_intf_84.fifo_rd_block = 0;
    assign fifo_intf_84.fifo_wr_block = 0;
    assign fifo_intf_84.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_84;
    csv_file_dump cstatus_csv_dumper_84;
    df_fifo_monitor fifo_monitor_84;
    df_fifo_intf fifo_intf_85(clock,reset);
    assign fifo_intf_85.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_3_U.if_empty_n;
    assign fifo_intf_85.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_3_U.if_full_n;
    assign fifo_intf_85.fifo_rd_block = 0;
    assign fifo_intf_85.fifo_wr_block = 0;
    assign fifo_intf_85.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_85;
    csv_file_dump cstatus_csv_dumper_85;
    df_fifo_monitor fifo_monitor_85;
    df_fifo_intf fifo_intf_86(clock,reset);
    assign fifo_intf_86.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_3_U.if_empty_n;
    assign fifo_intf_86.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_3_U.if_full_n;
    assign fifo_intf_86.fifo_rd_block = 0;
    assign fifo_intf_86.fifo_wr_block = 0;
    assign fifo_intf_86.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_86;
    csv_file_dump cstatus_csv_dumper_86;
    df_fifo_monitor fifo_monitor_86;
    df_fifo_intf fifo_intf_87(clock,reset);
    assign fifo_intf_87.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_3_U.if_empty_n;
    assign fifo_intf_87.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_3_U.if_full_n;
    assign fifo_intf_87.fifo_rd_block = 0;
    assign fifo_intf_87.fifo_wr_block = 0;
    assign fifo_intf_87.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_87;
    csv_file_dump cstatus_csv_dumper_87;
    df_fifo_monitor fifo_monitor_87;
    df_fifo_intf fifo_intf_88(clock,reset);
    assign fifo_intf_88.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_3_U.if_empty_n;
    assign fifo_intf_88.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_3_U.if_full_n;
    assign fifo_intf_88.fifo_rd_block = 0;
    assign fifo_intf_88.fifo_wr_block = 0;
    assign fifo_intf_88.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_88;
    csv_file_dump cstatus_csv_dumper_88;
    df_fifo_monitor fifo_monitor_88;
    df_fifo_intf fifo_intf_89(clock,reset);
    assign fifo_intf_89.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_3_U.if_empty_n;
    assign fifo_intf_89.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_3_U.if_full_n;
    assign fifo_intf_89.fifo_rd_block = 0;
    assign fifo_intf_89.fifo_wr_block = 0;
    assign fifo_intf_89.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_89;
    csv_file_dump cstatus_csv_dumper_89;
    df_fifo_monitor fifo_monitor_89;
    df_fifo_intf fifo_intf_90(clock,reset);
    assign fifo_intf_90.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_3_U.if_empty_n;
    assign fifo_intf_90.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_3_U.if_full_n;
    assign fifo_intf_90.fifo_rd_block = 0;
    assign fifo_intf_90.fifo_wr_block = 0;
    assign fifo_intf_90.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_90;
    csv_file_dump cstatus_csv_dumper_90;
    df_fifo_monitor fifo_monitor_90;
    df_fifo_intf fifo_intf_91(clock,reset);
    assign fifo_intf_91.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_3_U.if_empty_n;
    assign fifo_intf_91.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_3_U.if_full_n;
    assign fifo_intf_91.fifo_rd_block = 0;
    assign fifo_intf_91.fifo_wr_block = 0;
    assign fifo_intf_91.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_91;
    csv_file_dump cstatus_csv_dumper_91;
    df_fifo_monitor fifo_monitor_91;
    df_fifo_intf fifo_intf_92(clock,reset);
    assign fifo_intf_92.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_3_U.if_empty_n;
    assign fifo_intf_92.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_3_U.if_full_n;
    assign fifo_intf_92.fifo_rd_block = 0;
    assign fifo_intf_92.fifo_wr_block = 0;
    assign fifo_intf_92.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_92;
    csv_file_dump cstatus_csv_dumper_92;
    df_fifo_monitor fifo_monitor_92;
    df_fifo_intf fifo_intf_93(clock,reset);
    assign fifo_intf_93.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_3_U.if_empty_n;
    assign fifo_intf_93.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_3_U.if_full_n;
    assign fifo_intf_93.fifo_rd_block = 0;
    assign fifo_intf_93.fifo_wr_block = 0;
    assign fifo_intf_93.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_93;
    csv_file_dump cstatus_csv_dumper_93;
    df_fifo_monitor fifo_monitor_93;
    df_fifo_intf fifo_intf_94(clock,reset);
    assign fifo_intf_94.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_3_U.if_empty_n;
    assign fifo_intf_94.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_3_U.if_full_n;
    assign fifo_intf_94.fifo_rd_block = 0;
    assign fifo_intf_94.fifo_wr_block = 0;
    assign fifo_intf_94.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_94;
    csv_file_dump cstatus_csv_dumper_94;
    df_fifo_monitor fifo_monitor_94;
    df_fifo_intf fifo_intf_95(clock,reset);
    assign fifo_intf_95.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_3_U.if_empty_n;
    assign fifo_intf_95.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_3_U.if_full_n;
    assign fifo_intf_95.fifo_rd_block = 0;
    assign fifo_intf_95.fifo_wr_block = 0;
    assign fifo_intf_95.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_95;
    csv_file_dump cstatus_csv_dumper_95;
    df_fifo_monitor fifo_monitor_95;
    df_fifo_intf fifo_intf_96(clock,reset);
    assign fifo_intf_96.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_3_U.if_empty_n;
    assign fifo_intf_96.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_3_U.if_full_n;
    assign fifo_intf_96.fifo_rd_block = 0;
    assign fifo_intf_96.fifo_wr_block = 0;
    assign fifo_intf_96.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_96;
    csv_file_dump cstatus_csv_dumper_96;
    df_fifo_monitor fifo_monitor_96;
    df_fifo_intf fifo_intf_97(clock,reset);
    assign fifo_intf_97.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_3_U.if_empty_n;
    assign fifo_intf_97.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_3_U.if_full_n;
    assign fifo_intf_97.fifo_rd_block = 0;
    assign fifo_intf_97.fifo_wr_block = 0;
    assign fifo_intf_97.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_97;
    csv_file_dump cstatus_csv_dumper_97;
    df_fifo_monitor fifo_monitor_97;
    df_fifo_intf fifo_intf_98(clock,reset);
    assign fifo_intf_98.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_3_U.if_empty_n;
    assign fifo_intf_98.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_3_U.if_full_n;
    assign fifo_intf_98.fifo_rd_block = 0;
    assign fifo_intf_98.fifo_wr_block = 0;
    assign fifo_intf_98.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_98;
    csv_file_dump cstatus_csv_dumper_98;
    df_fifo_monitor fifo_monitor_98;
    df_fifo_intf fifo_intf_99(clock,reset);
    assign fifo_intf_99.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_3_U.if_empty_n;
    assign fifo_intf_99.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_3_U.if_full_n;
    assign fifo_intf_99.fifo_rd_block = 0;
    assign fifo_intf_99.fifo_wr_block = 0;
    assign fifo_intf_99.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_99;
    csv_file_dump cstatus_csv_dumper_99;
    df_fifo_monitor fifo_monitor_99;
    df_fifo_intf fifo_intf_100(clock,reset);
    assign fifo_intf_100.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_3_U.if_empty_n;
    assign fifo_intf_100.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_3_U.if_full_n;
    assign fifo_intf_100.fifo_rd_block = 0;
    assign fifo_intf_100.fifo_wr_block = 0;
    assign fifo_intf_100.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_100;
    csv_file_dump cstatus_csv_dumper_100;
    df_fifo_monitor fifo_monitor_100;
    df_fifo_intf fifo_intf_101(clock,reset);
    assign fifo_intf_101.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_3_U.if_empty_n;
    assign fifo_intf_101.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_3_U.if_full_n;
    assign fifo_intf_101.fifo_rd_block = 0;
    assign fifo_intf_101.fifo_wr_block = 0;
    assign fifo_intf_101.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_101;
    csv_file_dump cstatus_csv_dumper_101;
    df_fifo_monitor fifo_monitor_101;
    df_fifo_intf fifo_intf_102(clock,reset);
    assign fifo_intf_102.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_3_U.if_empty_n;
    assign fifo_intf_102.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_3_U.if_full_n;
    assign fifo_intf_102.fifo_rd_block = 0;
    assign fifo_intf_102.fifo_wr_block = 0;
    assign fifo_intf_102.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_102;
    csv_file_dump cstatus_csv_dumper_102;
    df_fifo_monitor fifo_monitor_102;
    df_fifo_intf fifo_intf_103(clock,reset);
    assign fifo_intf_103.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_4_U.if_empty_n;
    assign fifo_intf_103.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_4_U.if_full_n;
    assign fifo_intf_103.fifo_rd_block = 0;
    assign fifo_intf_103.fifo_wr_block = 0;
    assign fifo_intf_103.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_103;
    csv_file_dump cstatus_csv_dumper_103;
    df_fifo_monitor fifo_monitor_103;
    df_fifo_intf fifo_intf_104(clock,reset);
    assign fifo_intf_104.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_4_U.if_empty_n;
    assign fifo_intf_104.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_4_U.if_full_n;
    assign fifo_intf_104.fifo_rd_block = 0;
    assign fifo_intf_104.fifo_wr_block = 0;
    assign fifo_intf_104.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_104;
    csv_file_dump cstatus_csv_dumper_104;
    df_fifo_monitor fifo_monitor_104;
    df_fifo_intf fifo_intf_105(clock,reset);
    assign fifo_intf_105.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_4_U.if_empty_n;
    assign fifo_intf_105.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_4_U.if_full_n;
    assign fifo_intf_105.fifo_rd_block = 0;
    assign fifo_intf_105.fifo_wr_block = 0;
    assign fifo_intf_105.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_105;
    csv_file_dump cstatus_csv_dumper_105;
    df_fifo_monitor fifo_monitor_105;
    df_fifo_intf fifo_intf_106(clock,reset);
    assign fifo_intf_106.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_4_U.if_empty_n;
    assign fifo_intf_106.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_4_U.if_full_n;
    assign fifo_intf_106.fifo_rd_block = 0;
    assign fifo_intf_106.fifo_wr_block = 0;
    assign fifo_intf_106.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_106;
    csv_file_dump cstatus_csv_dumper_106;
    df_fifo_monitor fifo_monitor_106;
    df_fifo_intf fifo_intf_107(clock,reset);
    assign fifo_intf_107.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_4_U.if_empty_n;
    assign fifo_intf_107.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_4_U.if_full_n;
    assign fifo_intf_107.fifo_rd_block = 0;
    assign fifo_intf_107.fifo_wr_block = 0;
    assign fifo_intf_107.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_107;
    csv_file_dump cstatus_csv_dumper_107;
    df_fifo_monitor fifo_monitor_107;
    df_fifo_intf fifo_intf_108(clock,reset);
    assign fifo_intf_108.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_4_U.if_empty_n;
    assign fifo_intf_108.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_4_U.if_full_n;
    assign fifo_intf_108.fifo_rd_block = 0;
    assign fifo_intf_108.fifo_wr_block = 0;
    assign fifo_intf_108.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_108;
    csv_file_dump cstatus_csv_dumper_108;
    df_fifo_monitor fifo_monitor_108;
    df_fifo_intf fifo_intf_109(clock,reset);
    assign fifo_intf_109.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_4_U.if_empty_n;
    assign fifo_intf_109.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_4_U.if_full_n;
    assign fifo_intf_109.fifo_rd_block = 0;
    assign fifo_intf_109.fifo_wr_block = 0;
    assign fifo_intf_109.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_109;
    csv_file_dump cstatus_csv_dumper_109;
    df_fifo_monitor fifo_monitor_109;
    df_fifo_intf fifo_intf_110(clock,reset);
    assign fifo_intf_110.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_4_U.if_empty_n;
    assign fifo_intf_110.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_4_U.if_full_n;
    assign fifo_intf_110.fifo_rd_block = 0;
    assign fifo_intf_110.fifo_wr_block = 0;
    assign fifo_intf_110.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_110;
    csv_file_dump cstatus_csv_dumper_110;
    df_fifo_monitor fifo_monitor_110;
    df_fifo_intf fifo_intf_111(clock,reset);
    assign fifo_intf_111.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_4_U.if_empty_n;
    assign fifo_intf_111.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_4_U.if_full_n;
    assign fifo_intf_111.fifo_rd_block = 0;
    assign fifo_intf_111.fifo_wr_block = 0;
    assign fifo_intf_111.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_111;
    csv_file_dump cstatus_csv_dumper_111;
    df_fifo_monitor fifo_monitor_111;
    df_fifo_intf fifo_intf_112(clock,reset);
    assign fifo_intf_112.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_4_U.if_empty_n;
    assign fifo_intf_112.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_4_U.if_full_n;
    assign fifo_intf_112.fifo_rd_block = 0;
    assign fifo_intf_112.fifo_wr_block = 0;
    assign fifo_intf_112.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_112;
    csv_file_dump cstatus_csv_dumper_112;
    df_fifo_monitor fifo_monitor_112;
    df_fifo_intf fifo_intf_113(clock,reset);
    assign fifo_intf_113.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_4_U.if_empty_n;
    assign fifo_intf_113.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_4_U.if_full_n;
    assign fifo_intf_113.fifo_rd_block = 0;
    assign fifo_intf_113.fifo_wr_block = 0;
    assign fifo_intf_113.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_113;
    csv_file_dump cstatus_csv_dumper_113;
    df_fifo_monitor fifo_monitor_113;
    df_fifo_intf fifo_intf_114(clock,reset);
    assign fifo_intf_114.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_4_U.if_empty_n;
    assign fifo_intf_114.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_4_U.if_full_n;
    assign fifo_intf_114.fifo_rd_block = 0;
    assign fifo_intf_114.fifo_wr_block = 0;
    assign fifo_intf_114.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_114;
    csv_file_dump cstatus_csv_dumper_114;
    df_fifo_monitor fifo_monitor_114;
    df_fifo_intf fifo_intf_115(clock,reset);
    assign fifo_intf_115.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_4_U.if_empty_n;
    assign fifo_intf_115.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_4_U.if_full_n;
    assign fifo_intf_115.fifo_rd_block = 0;
    assign fifo_intf_115.fifo_wr_block = 0;
    assign fifo_intf_115.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_115;
    csv_file_dump cstatus_csv_dumper_115;
    df_fifo_monitor fifo_monitor_115;
    df_fifo_intf fifo_intf_116(clock,reset);
    assign fifo_intf_116.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_4_U.if_empty_n;
    assign fifo_intf_116.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_4_U.if_full_n;
    assign fifo_intf_116.fifo_rd_block = 0;
    assign fifo_intf_116.fifo_wr_block = 0;
    assign fifo_intf_116.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_116;
    csv_file_dump cstatus_csv_dumper_116;
    df_fifo_monitor fifo_monitor_116;
    df_fifo_intf fifo_intf_117(clock,reset);
    assign fifo_intf_117.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_4_U.if_empty_n;
    assign fifo_intf_117.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_4_U.if_full_n;
    assign fifo_intf_117.fifo_rd_block = 0;
    assign fifo_intf_117.fifo_wr_block = 0;
    assign fifo_intf_117.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_117;
    csv_file_dump cstatus_csv_dumper_117;
    df_fifo_monitor fifo_monitor_117;
    df_fifo_intf fifo_intf_118(clock,reset);
    assign fifo_intf_118.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_4_U.if_empty_n;
    assign fifo_intf_118.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_4_U.if_full_n;
    assign fifo_intf_118.fifo_rd_block = 0;
    assign fifo_intf_118.fifo_wr_block = 0;
    assign fifo_intf_118.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_118;
    csv_file_dump cstatus_csv_dumper_118;
    df_fifo_monitor fifo_monitor_118;
    df_fifo_intf fifo_intf_119(clock,reset);
    assign fifo_intf_119.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_4_U.if_empty_n;
    assign fifo_intf_119.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_4_U.if_full_n;
    assign fifo_intf_119.fifo_rd_block = 0;
    assign fifo_intf_119.fifo_wr_block = 0;
    assign fifo_intf_119.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_119;
    csv_file_dump cstatus_csv_dumper_119;
    df_fifo_monitor fifo_monitor_119;
    df_fifo_intf fifo_intf_120(clock,reset);
    assign fifo_intf_120.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_4_U.if_empty_n;
    assign fifo_intf_120.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_4_U.if_full_n;
    assign fifo_intf_120.fifo_rd_block = 0;
    assign fifo_intf_120.fifo_wr_block = 0;
    assign fifo_intf_120.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_120;
    csv_file_dump cstatus_csv_dumper_120;
    df_fifo_monitor fifo_monitor_120;
    df_fifo_intf fifo_intf_121(clock,reset);
    assign fifo_intf_121.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_4_U.if_empty_n;
    assign fifo_intf_121.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_4_U.if_full_n;
    assign fifo_intf_121.fifo_rd_block = 0;
    assign fifo_intf_121.fifo_wr_block = 0;
    assign fifo_intf_121.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_121;
    csv_file_dump cstatus_csv_dumper_121;
    df_fifo_monitor fifo_monitor_121;
    df_fifo_intf fifo_intf_122(clock,reset);
    assign fifo_intf_122.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_4_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_4_U.if_empty_n;
    assign fifo_intf_122.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_4_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_4_U.if_full_n;
    assign fifo_intf_122.fifo_rd_block = 0;
    assign fifo_intf_122.fifo_wr_block = 0;
    assign fifo_intf_122.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_122;
    csv_file_dump cstatus_csv_dumper_122;
    df_fifo_monitor fifo_monitor_122;
    df_fifo_intf fifo_intf_123(clock,reset);
    assign fifo_intf_123.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_5_U.if_empty_n;
    assign fifo_intf_123.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_5_U.if_full_n;
    assign fifo_intf_123.fifo_rd_block = 0;
    assign fifo_intf_123.fifo_wr_block = 0;
    assign fifo_intf_123.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_123;
    csv_file_dump cstatus_csv_dumper_123;
    df_fifo_monitor fifo_monitor_123;
    df_fifo_intf fifo_intf_124(clock,reset);
    assign fifo_intf_124.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_5_U.if_empty_n;
    assign fifo_intf_124.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_5_U.if_full_n;
    assign fifo_intf_124.fifo_rd_block = 0;
    assign fifo_intf_124.fifo_wr_block = 0;
    assign fifo_intf_124.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_124;
    csv_file_dump cstatus_csv_dumper_124;
    df_fifo_monitor fifo_monitor_124;
    df_fifo_intf fifo_intf_125(clock,reset);
    assign fifo_intf_125.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_5_U.if_empty_n;
    assign fifo_intf_125.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_5_U.if_full_n;
    assign fifo_intf_125.fifo_rd_block = 0;
    assign fifo_intf_125.fifo_wr_block = 0;
    assign fifo_intf_125.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_125;
    csv_file_dump cstatus_csv_dumper_125;
    df_fifo_monitor fifo_monitor_125;
    df_fifo_intf fifo_intf_126(clock,reset);
    assign fifo_intf_126.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_5_U.if_empty_n;
    assign fifo_intf_126.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_5_U.if_full_n;
    assign fifo_intf_126.fifo_rd_block = 0;
    assign fifo_intf_126.fifo_wr_block = 0;
    assign fifo_intf_126.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_126;
    csv_file_dump cstatus_csv_dumper_126;
    df_fifo_monitor fifo_monitor_126;
    df_fifo_intf fifo_intf_127(clock,reset);
    assign fifo_intf_127.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_5_U.if_empty_n;
    assign fifo_intf_127.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_5_U.if_full_n;
    assign fifo_intf_127.fifo_rd_block = 0;
    assign fifo_intf_127.fifo_wr_block = 0;
    assign fifo_intf_127.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_127;
    csv_file_dump cstatus_csv_dumper_127;
    df_fifo_monitor fifo_monitor_127;
    df_fifo_intf fifo_intf_128(clock,reset);
    assign fifo_intf_128.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_5_U.if_empty_n;
    assign fifo_intf_128.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_5_U.if_full_n;
    assign fifo_intf_128.fifo_rd_block = 0;
    assign fifo_intf_128.fifo_wr_block = 0;
    assign fifo_intf_128.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_128;
    csv_file_dump cstatus_csv_dumper_128;
    df_fifo_monitor fifo_monitor_128;
    df_fifo_intf fifo_intf_129(clock,reset);
    assign fifo_intf_129.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_5_U.if_empty_n;
    assign fifo_intf_129.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_5_U.if_full_n;
    assign fifo_intf_129.fifo_rd_block = 0;
    assign fifo_intf_129.fifo_wr_block = 0;
    assign fifo_intf_129.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_129;
    csv_file_dump cstatus_csv_dumper_129;
    df_fifo_monitor fifo_monitor_129;
    df_fifo_intf fifo_intf_130(clock,reset);
    assign fifo_intf_130.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_5_U.if_empty_n;
    assign fifo_intf_130.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_5_U.if_full_n;
    assign fifo_intf_130.fifo_rd_block = 0;
    assign fifo_intf_130.fifo_wr_block = 0;
    assign fifo_intf_130.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_130;
    csv_file_dump cstatus_csv_dumper_130;
    df_fifo_monitor fifo_monitor_130;
    df_fifo_intf fifo_intf_131(clock,reset);
    assign fifo_intf_131.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_5_U.if_empty_n;
    assign fifo_intf_131.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_5_U.if_full_n;
    assign fifo_intf_131.fifo_rd_block = 0;
    assign fifo_intf_131.fifo_wr_block = 0;
    assign fifo_intf_131.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_131;
    csv_file_dump cstatus_csv_dumper_131;
    df_fifo_monitor fifo_monitor_131;
    df_fifo_intf fifo_intf_132(clock,reset);
    assign fifo_intf_132.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_5_U.if_empty_n;
    assign fifo_intf_132.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_5_U.if_full_n;
    assign fifo_intf_132.fifo_rd_block = 0;
    assign fifo_intf_132.fifo_wr_block = 0;
    assign fifo_intf_132.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_132;
    csv_file_dump cstatus_csv_dumper_132;
    df_fifo_monitor fifo_monitor_132;
    df_fifo_intf fifo_intf_133(clock,reset);
    assign fifo_intf_133.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_5_U.if_empty_n;
    assign fifo_intf_133.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_5_U.if_full_n;
    assign fifo_intf_133.fifo_rd_block = 0;
    assign fifo_intf_133.fifo_wr_block = 0;
    assign fifo_intf_133.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_133;
    csv_file_dump cstatus_csv_dumper_133;
    df_fifo_monitor fifo_monitor_133;
    df_fifo_intf fifo_intf_134(clock,reset);
    assign fifo_intf_134.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_5_U.if_empty_n;
    assign fifo_intf_134.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_5_U.if_full_n;
    assign fifo_intf_134.fifo_rd_block = 0;
    assign fifo_intf_134.fifo_wr_block = 0;
    assign fifo_intf_134.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_134;
    csv_file_dump cstatus_csv_dumper_134;
    df_fifo_monitor fifo_monitor_134;
    df_fifo_intf fifo_intf_135(clock,reset);
    assign fifo_intf_135.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_5_U.if_empty_n;
    assign fifo_intf_135.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_5_U.if_full_n;
    assign fifo_intf_135.fifo_rd_block = 0;
    assign fifo_intf_135.fifo_wr_block = 0;
    assign fifo_intf_135.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_135;
    csv_file_dump cstatus_csv_dumper_135;
    df_fifo_monitor fifo_monitor_135;
    df_fifo_intf fifo_intf_136(clock,reset);
    assign fifo_intf_136.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_5_U.if_empty_n;
    assign fifo_intf_136.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_5_U.if_full_n;
    assign fifo_intf_136.fifo_rd_block = 0;
    assign fifo_intf_136.fifo_wr_block = 0;
    assign fifo_intf_136.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_136;
    csv_file_dump cstatus_csv_dumper_136;
    df_fifo_monitor fifo_monitor_136;
    df_fifo_intf fifo_intf_137(clock,reset);
    assign fifo_intf_137.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_5_U.if_empty_n;
    assign fifo_intf_137.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_5_U.if_full_n;
    assign fifo_intf_137.fifo_rd_block = 0;
    assign fifo_intf_137.fifo_wr_block = 0;
    assign fifo_intf_137.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_137;
    csv_file_dump cstatus_csv_dumper_137;
    df_fifo_monitor fifo_monitor_137;
    df_fifo_intf fifo_intf_138(clock,reset);
    assign fifo_intf_138.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_5_U.if_empty_n;
    assign fifo_intf_138.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_5_U.if_full_n;
    assign fifo_intf_138.fifo_rd_block = 0;
    assign fifo_intf_138.fifo_wr_block = 0;
    assign fifo_intf_138.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_138;
    csv_file_dump cstatus_csv_dumper_138;
    df_fifo_monitor fifo_monitor_138;
    df_fifo_intf fifo_intf_139(clock,reset);
    assign fifo_intf_139.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_5_U.if_empty_n;
    assign fifo_intf_139.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_5_U.if_full_n;
    assign fifo_intf_139.fifo_rd_block = 0;
    assign fifo_intf_139.fifo_wr_block = 0;
    assign fifo_intf_139.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_139;
    csv_file_dump cstatus_csv_dumper_139;
    df_fifo_monitor fifo_monitor_139;
    df_fifo_intf fifo_intf_140(clock,reset);
    assign fifo_intf_140.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_5_U.if_empty_n;
    assign fifo_intf_140.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_5_U.if_full_n;
    assign fifo_intf_140.fifo_rd_block = 0;
    assign fifo_intf_140.fifo_wr_block = 0;
    assign fifo_intf_140.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_140;
    csv_file_dump cstatus_csv_dumper_140;
    df_fifo_monitor fifo_monitor_140;
    df_fifo_intf fifo_intf_141(clock,reset);
    assign fifo_intf_141.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_5_U.if_empty_n;
    assign fifo_intf_141.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_5_U.if_full_n;
    assign fifo_intf_141.fifo_rd_block = 0;
    assign fifo_intf_141.fifo_wr_block = 0;
    assign fifo_intf_141.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_141;
    csv_file_dump cstatus_csv_dumper_141;
    df_fifo_monitor fifo_monitor_141;
    df_fifo_intf fifo_intf_142(clock,reset);
    assign fifo_intf_142.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_5_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_5_U.if_empty_n;
    assign fifo_intf_142.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_5_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_5_U.if_full_n;
    assign fifo_intf_142.fifo_rd_block = 0;
    assign fifo_intf_142.fifo_wr_block = 0;
    assign fifo_intf_142.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_142;
    csv_file_dump cstatus_csv_dumper_142;
    df_fifo_monitor fifo_monitor_142;
    df_fifo_intf fifo_intf_143(clock,reset);
    assign fifo_intf_143.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_6_U.if_empty_n;
    assign fifo_intf_143.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_6_U.if_full_n;
    assign fifo_intf_143.fifo_rd_block = 0;
    assign fifo_intf_143.fifo_wr_block = 0;
    assign fifo_intf_143.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_143;
    csv_file_dump cstatus_csv_dumper_143;
    df_fifo_monitor fifo_monitor_143;
    df_fifo_intf fifo_intf_144(clock,reset);
    assign fifo_intf_144.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_6_U.if_empty_n;
    assign fifo_intf_144.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_6_U.if_full_n;
    assign fifo_intf_144.fifo_rd_block = 0;
    assign fifo_intf_144.fifo_wr_block = 0;
    assign fifo_intf_144.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_144;
    csv_file_dump cstatus_csv_dumper_144;
    df_fifo_monitor fifo_monitor_144;
    df_fifo_intf fifo_intf_145(clock,reset);
    assign fifo_intf_145.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_6_U.if_empty_n;
    assign fifo_intf_145.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_6_U.if_full_n;
    assign fifo_intf_145.fifo_rd_block = 0;
    assign fifo_intf_145.fifo_wr_block = 0;
    assign fifo_intf_145.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_145;
    csv_file_dump cstatus_csv_dumper_145;
    df_fifo_monitor fifo_monitor_145;
    df_fifo_intf fifo_intf_146(clock,reset);
    assign fifo_intf_146.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_6_U.if_empty_n;
    assign fifo_intf_146.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_6_U.if_full_n;
    assign fifo_intf_146.fifo_rd_block = 0;
    assign fifo_intf_146.fifo_wr_block = 0;
    assign fifo_intf_146.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_146;
    csv_file_dump cstatus_csv_dumper_146;
    df_fifo_monitor fifo_monitor_146;
    df_fifo_intf fifo_intf_147(clock,reset);
    assign fifo_intf_147.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_6_U.if_empty_n;
    assign fifo_intf_147.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_6_U.if_full_n;
    assign fifo_intf_147.fifo_rd_block = 0;
    assign fifo_intf_147.fifo_wr_block = 0;
    assign fifo_intf_147.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_147;
    csv_file_dump cstatus_csv_dumper_147;
    df_fifo_monitor fifo_monitor_147;
    df_fifo_intf fifo_intf_148(clock,reset);
    assign fifo_intf_148.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_6_U.if_empty_n;
    assign fifo_intf_148.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_6_U.if_full_n;
    assign fifo_intf_148.fifo_rd_block = 0;
    assign fifo_intf_148.fifo_wr_block = 0;
    assign fifo_intf_148.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_148;
    csv_file_dump cstatus_csv_dumper_148;
    df_fifo_monitor fifo_monitor_148;
    df_fifo_intf fifo_intf_149(clock,reset);
    assign fifo_intf_149.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_6_U.if_empty_n;
    assign fifo_intf_149.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_6_U.if_full_n;
    assign fifo_intf_149.fifo_rd_block = 0;
    assign fifo_intf_149.fifo_wr_block = 0;
    assign fifo_intf_149.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_149;
    csv_file_dump cstatus_csv_dumper_149;
    df_fifo_monitor fifo_monitor_149;
    df_fifo_intf fifo_intf_150(clock,reset);
    assign fifo_intf_150.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_6_U.if_empty_n;
    assign fifo_intf_150.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_6_U.if_full_n;
    assign fifo_intf_150.fifo_rd_block = 0;
    assign fifo_intf_150.fifo_wr_block = 0;
    assign fifo_intf_150.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_150;
    csv_file_dump cstatus_csv_dumper_150;
    df_fifo_monitor fifo_monitor_150;
    df_fifo_intf fifo_intf_151(clock,reset);
    assign fifo_intf_151.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_6_U.if_empty_n;
    assign fifo_intf_151.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_6_U.if_full_n;
    assign fifo_intf_151.fifo_rd_block = 0;
    assign fifo_intf_151.fifo_wr_block = 0;
    assign fifo_intf_151.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_151;
    csv_file_dump cstatus_csv_dumper_151;
    df_fifo_monitor fifo_monitor_151;
    df_fifo_intf fifo_intf_152(clock,reset);
    assign fifo_intf_152.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_6_U.if_empty_n;
    assign fifo_intf_152.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_6_U.if_full_n;
    assign fifo_intf_152.fifo_rd_block = 0;
    assign fifo_intf_152.fifo_wr_block = 0;
    assign fifo_intf_152.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_152;
    csv_file_dump cstatus_csv_dumper_152;
    df_fifo_monitor fifo_monitor_152;
    df_fifo_intf fifo_intf_153(clock,reset);
    assign fifo_intf_153.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_6_U.if_empty_n;
    assign fifo_intf_153.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_6_U.if_full_n;
    assign fifo_intf_153.fifo_rd_block = 0;
    assign fifo_intf_153.fifo_wr_block = 0;
    assign fifo_intf_153.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_153;
    csv_file_dump cstatus_csv_dumper_153;
    df_fifo_monitor fifo_monitor_153;
    df_fifo_intf fifo_intf_154(clock,reset);
    assign fifo_intf_154.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_6_U.if_empty_n;
    assign fifo_intf_154.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_6_U.if_full_n;
    assign fifo_intf_154.fifo_rd_block = 0;
    assign fifo_intf_154.fifo_wr_block = 0;
    assign fifo_intf_154.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_154;
    csv_file_dump cstatus_csv_dumper_154;
    df_fifo_monitor fifo_monitor_154;
    df_fifo_intf fifo_intf_155(clock,reset);
    assign fifo_intf_155.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_6_U.if_empty_n;
    assign fifo_intf_155.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_6_U.if_full_n;
    assign fifo_intf_155.fifo_rd_block = 0;
    assign fifo_intf_155.fifo_wr_block = 0;
    assign fifo_intf_155.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_155;
    csv_file_dump cstatus_csv_dumper_155;
    df_fifo_monitor fifo_monitor_155;
    df_fifo_intf fifo_intf_156(clock,reset);
    assign fifo_intf_156.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_6_U.if_empty_n;
    assign fifo_intf_156.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_6_U.if_full_n;
    assign fifo_intf_156.fifo_rd_block = 0;
    assign fifo_intf_156.fifo_wr_block = 0;
    assign fifo_intf_156.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_156;
    csv_file_dump cstatus_csv_dumper_156;
    df_fifo_monitor fifo_monitor_156;
    df_fifo_intf fifo_intf_157(clock,reset);
    assign fifo_intf_157.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_6_U.if_empty_n;
    assign fifo_intf_157.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_6_U.if_full_n;
    assign fifo_intf_157.fifo_rd_block = 0;
    assign fifo_intf_157.fifo_wr_block = 0;
    assign fifo_intf_157.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_157;
    csv_file_dump cstatus_csv_dumper_157;
    df_fifo_monitor fifo_monitor_157;
    df_fifo_intf fifo_intf_158(clock,reset);
    assign fifo_intf_158.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_6_U.if_empty_n;
    assign fifo_intf_158.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_6_U.if_full_n;
    assign fifo_intf_158.fifo_rd_block = 0;
    assign fifo_intf_158.fifo_wr_block = 0;
    assign fifo_intf_158.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_158;
    csv_file_dump cstatus_csv_dumper_158;
    df_fifo_monitor fifo_monitor_158;
    df_fifo_intf fifo_intf_159(clock,reset);
    assign fifo_intf_159.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_6_U.if_empty_n;
    assign fifo_intf_159.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_6_U.if_full_n;
    assign fifo_intf_159.fifo_rd_block = 0;
    assign fifo_intf_159.fifo_wr_block = 0;
    assign fifo_intf_159.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_159;
    csv_file_dump cstatus_csv_dumper_159;
    df_fifo_monitor fifo_monitor_159;
    df_fifo_intf fifo_intf_160(clock,reset);
    assign fifo_intf_160.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_6_U.if_empty_n;
    assign fifo_intf_160.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_6_U.if_full_n;
    assign fifo_intf_160.fifo_rd_block = 0;
    assign fifo_intf_160.fifo_wr_block = 0;
    assign fifo_intf_160.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_160;
    csv_file_dump cstatus_csv_dumper_160;
    df_fifo_monitor fifo_monitor_160;
    df_fifo_intf fifo_intf_161(clock,reset);
    assign fifo_intf_161.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_6_U.if_empty_n;
    assign fifo_intf_161.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_6_U.if_full_n;
    assign fifo_intf_161.fifo_rd_block = 0;
    assign fifo_intf_161.fifo_wr_block = 0;
    assign fifo_intf_161.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_161;
    csv_file_dump cstatus_csv_dumper_161;
    df_fifo_monitor fifo_monitor_161;
    df_fifo_intf fifo_intf_162(clock,reset);
    assign fifo_intf_162.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_6_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_6_U.if_empty_n;
    assign fifo_intf_162.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_6_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_6_U.if_full_n;
    assign fifo_intf_162.fifo_rd_block = 0;
    assign fifo_intf_162.fifo_wr_block = 0;
    assign fifo_intf_162.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_162;
    csv_file_dump cstatus_csv_dumper_162;
    df_fifo_monitor fifo_monitor_162;
    df_fifo_intf fifo_intf_163(clock,reset);
    assign fifo_intf_163.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_7_U.if_empty_n;
    assign fifo_intf_163.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_7_U.if_full_n;
    assign fifo_intf_163.fifo_rd_block = 0;
    assign fifo_intf_163.fifo_wr_block = 0;
    assign fifo_intf_163.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_163;
    csv_file_dump cstatus_csv_dumper_163;
    df_fifo_monitor fifo_monitor_163;
    df_fifo_intf fifo_intf_164(clock,reset);
    assign fifo_intf_164.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_7_U.if_empty_n;
    assign fifo_intf_164.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_7_U.if_full_n;
    assign fifo_intf_164.fifo_rd_block = 0;
    assign fifo_intf_164.fifo_wr_block = 0;
    assign fifo_intf_164.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_164;
    csv_file_dump cstatus_csv_dumper_164;
    df_fifo_monitor fifo_monitor_164;
    df_fifo_intf fifo_intf_165(clock,reset);
    assign fifo_intf_165.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_7_U.if_empty_n;
    assign fifo_intf_165.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_7_U.if_full_n;
    assign fifo_intf_165.fifo_rd_block = 0;
    assign fifo_intf_165.fifo_wr_block = 0;
    assign fifo_intf_165.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_165;
    csv_file_dump cstatus_csv_dumper_165;
    df_fifo_monitor fifo_monitor_165;
    df_fifo_intf fifo_intf_166(clock,reset);
    assign fifo_intf_166.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_7_U.if_empty_n;
    assign fifo_intf_166.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_7_U.if_full_n;
    assign fifo_intf_166.fifo_rd_block = 0;
    assign fifo_intf_166.fifo_wr_block = 0;
    assign fifo_intf_166.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_166;
    csv_file_dump cstatus_csv_dumper_166;
    df_fifo_monitor fifo_monitor_166;
    df_fifo_intf fifo_intf_167(clock,reset);
    assign fifo_intf_167.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_7_U.if_empty_n;
    assign fifo_intf_167.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_7_U.if_full_n;
    assign fifo_intf_167.fifo_rd_block = 0;
    assign fifo_intf_167.fifo_wr_block = 0;
    assign fifo_intf_167.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_167;
    csv_file_dump cstatus_csv_dumper_167;
    df_fifo_monitor fifo_monitor_167;
    df_fifo_intf fifo_intf_168(clock,reset);
    assign fifo_intf_168.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_7_U.if_empty_n;
    assign fifo_intf_168.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_7_U.if_full_n;
    assign fifo_intf_168.fifo_rd_block = 0;
    assign fifo_intf_168.fifo_wr_block = 0;
    assign fifo_intf_168.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_168;
    csv_file_dump cstatus_csv_dumper_168;
    df_fifo_monitor fifo_monitor_168;
    df_fifo_intf fifo_intf_169(clock,reset);
    assign fifo_intf_169.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_7_U.if_empty_n;
    assign fifo_intf_169.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_7_U.if_full_n;
    assign fifo_intf_169.fifo_rd_block = 0;
    assign fifo_intf_169.fifo_wr_block = 0;
    assign fifo_intf_169.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_169;
    csv_file_dump cstatus_csv_dumper_169;
    df_fifo_monitor fifo_monitor_169;
    df_fifo_intf fifo_intf_170(clock,reset);
    assign fifo_intf_170.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_7_U.if_empty_n;
    assign fifo_intf_170.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_7_U.if_full_n;
    assign fifo_intf_170.fifo_rd_block = 0;
    assign fifo_intf_170.fifo_wr_block = 0;
    assign fifo_intf_170.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_170;
    csv_file_dump cstatus_csv_dumper_170;
    df_fifo_monitor fifo_monitor_170;
    df_fifo_intf fifo_intf_171(clock,reset);
    assign fifo_intf_171.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_7_U.if_empty_n;
    assign fifo_intf_171.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_7_U.if_full_n;
    assign fifo_intf_171.fifo_rd_block = 0;
    assign fifo_intf_171.fifo_wr_block = 0;
    assign fifo_intf_171.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_171;
    csv_file_dump cstatus_csv_dumper_171;
    df_fifo_monitor fifo_monitor_171;
    df_fifo_intf fifo_intf_172(clock,reset);
    assign fifo_intf_172.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_7_U.if_empty_n;
    assign fifo_intf_172.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_7_U.if_full_n;
    assign fifo_intf_172.fifo_rd_block = 0;
    assign fifo_intf_172.fifo_wr_block = 0;
    assign fifo_intf_172.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_172;
    csv_file_dump cstatus_csv_dumper_172;
    df_fifo_monitor fifo_monitor_172;
    df_fifo_intf fifo_intf_173(clock,reset);
    assign fifo_intf_173.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_7_U.if_empty_n;
    assign fifo_intf_173.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_7_U.if_full_n;
    assign fifo_intf_173.fifo_rd_block = 0;
    assign fifo_intf_173.fifo_wr_block = 0;
    assign fifo_intf_173.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_173;
    csv_file_dump cstatus_csv_dumper_173;
    df_fifo_monitor fifo_monitor_173;
    df_fifo_intf fifo_intf_174(clock,reset);
    assign fifo_intf_174.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_7_U.if_empty_n;
    assign fifo_intf_174.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_7_U.if_full_n;
    assign fifo_intf_174.fifo_rd_block = 0;
    assign fifo_intf_174.fifo_wr_block = 0;
    assign fifo_intf_174.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_174;
    csv_file_dump cstatus_csv_dumper_174;
    df_fifo_monitor fifo_monitor_174;
    df_fifo_intf fifo_intf_175(clock,reset);
    assign fifo_intf_175.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_7_U.if_empty_n;
    assign fifo_intf_175.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_7_U.if_full_n;
    assign fifo_intf_175.fifo_rd_block = 0;
    assign fifo_intf_175.fifo_wr_block = 0;
    assign fifo_intf_175.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_175;
    csv_file_dump cstatus_csv_dumper_175;
    df_fifo_monitor fifo_monitor_175;
    df_fifo_intf fifo_intf_176(clock,reset);
    assign fifo_intf_176.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_7_U.if_empty_n;
    assign fifo_intf_176.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_7_U.if_full_n;
    assign fifo_intf_176.fifo_rd_block = 0;
    assign fifo_intf_176.fifo_wr_block = 0;
    assign fifo_intf_176.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_176;
    csv_file_dump cstatus_csv_dumper_176;
    df_fifo_monitor fifo_monitor_176;
    df_fifo_intf fifo_intf_177(clock,reset);
    assign fifo_intf_177.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_7_U.if_empty_n;
    assign fifo_intf_177.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_7_U.if_full_n;
    assign fifo_intf_177.fifo_rd_block = 0;
    assign fifo_intf_177.fifo_wr_block = 0;
    assign fifo_intf_177.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_177;
    csv_file_dump cstatus_csv_dumper_177;
    df_fifo_monitor fifo_monitor_177;
    df_fifo_intf fifo_intf_178(clock,reset);
    assign fifo_intf_178.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_7_U.if_empty_n;
    assign fifo_intf_178.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_7_U.if_full_n;
    assign fifo_intf_178.fifo_rd_block = 0;
    assign fifo_intf_178.fifo_wr_block = 0;
    assign fifo_intf_178.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_178;
    csv_file_dump cstatus_csv_dumper_178;
    df_fifo_monitor fifo_monitor_178;
    df_fifo_intf fifo_intf_179(clock,reset);
    assign fifo_intf_179.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_7_U.if_empty_n;
    assign fifo_intf_179.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_7_U.if_full_n;
    assign fifo_intf_179.fifo_rd_block = 0;
    assign fifo_intf_179.fifo_wr_block = 0;
    assign fifo_intf_179.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_179;
    csv_file_dump cstatus_csv_dumper_179;
    df_fifo_monitor fifo_monitor_179;
    df_fifo_intf fifo_intf_180(clock,reset);
    assign fifo_intf_180.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_7_U.if_empty_n;
    assign fifo_intf_180.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_7_U.if_full_n;
    assign fifo_intf_180.fifo_rd_block = 0;
    assign fifo_intf_180.fifo_wr_block = 0;
    assign fifo_intf_180.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_180;
    csv_file_dump cstatus_csv_dumper_180;
    df_fifo_monitor fifo_monitor_180;
    df_fifo_intf fifo_intf_181(clock,reset);
    assign fifo_intf_181.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_7_U.if_empty_n;
    assign fifo_intf_181.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_7_U.if_full_n;
    assign fifo_intf_181.fifo_rd_block = 0;
    assign fifo_intf_181.fifo_wr_block = 0;
    assign fifo_intf_181.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_181;
    csv_file_dump cstatus_csv_dumper_181;
    df_fifo_monitor fifo_monitor_181;
    df_fifo_intf fifo_intf_182(clock,reset);
    assign fifo_intf_182.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_7_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_7_U.if_empty_n;
    assign fifo_intf_182.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_7_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_7_U.if_full_n;
    assign fifo_intf_182.fifo_rd_block = 0;
    assign fifo_intf_182.fifo_wr_block = 0;
    assign fifo_intf_182.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_182;
    csv_file_dump cstatus_csv_dumper_182;
    df_fifo_monitor fifo_monitor_182;
    df_fifo_intf fifo_intf_183(clock,reset);
    assign fifo_intf_183.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_8_U.if_empty_n;
    assign fifo_intf_183.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_8_U.if_full_n;
    assign fifo_intf_183.fifo_rd_block = 0;
    assign fifo_intf_183.fifo_wr_block = 0;
    assign fifo_intf_183.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_183;
    csv_file_dump cstatus_csv_dumper_183;
    df_fifo_monitor fifo_monitor_183;
    df_fifo_intf fifo_intf_184(clock,reset);
    assign fifo_intf_184.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_8_U.if_empty_n;
    assign fifo_intf_184.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_8_U.if_full_n;
    assign fifo_intf_184.fifo_rd_block = 0;
    assign fifo_intf_184.fifo_wr_block = 0;
    assign fifo_intf_184.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_184;
    csv_file_dump cstatus_csv_dumper_184;
    df_fifo_monitor fifo_monitor_184;
    df_fifo_intf fifo_intf_185(clock,reset);
    assign fifo_intf_185.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_8_U.if_empty_n;
    assign fifo_intf_185.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_8_U.if_full_n;
    assign fifo_intf_185.fifo_rd_block = 0;
    assign fifo_intf_185.fifo_wr_block = 0;
    assign fifo_intf_185.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_185;
    csv_file_dump cstatus_csv_dumper_185;
    df_fifo_monitor fifo_monitor_185;
    df_fifo_intf fifo_intf_186(clock,reset);
    assign fifo_intf_186.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_8_U.if_empty_n;
    assign fifo_intf_186.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_8_U.if_full_n;
    assign fifo_intf_186.fifo_rd_block = 0;
    assign fifo_intf_186.fifo_wr_block = 0;
    assign fifo_intf_186.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_186;
    csv_file_dump cstatus_csv_dumper_186;
    df_fifo_monitor fifo_monitor_186;
    df_fifo_intf fifo_intf_187(clock,reset);
    assign fifo_intf_187.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_8_U.if_empty_n;
    assign fifo_intf_187.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_8_U.if_full_n;
    assign fifo_intf_187.fifo_rd_block = 0;
    assign fifo_intf_187.fifo_wr_block = 0;
    assign fifo_intf_187.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_187;
    csv_file_dump cstatus_csv_dumper_187;
    df_fifo_monitor fifo_monitor_187;
    df_fifo_intf fifo_intf_188(clock,reset);
    assign fifo_intf_188.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_8_U.if_empty_n;
    assign fifo_intf_188.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_8_U.if_full_n;
    assign fifo_intf_188.fifo_rd_block = 0;
    assign fifo_intf_188.fifo_wr_block = 0;
    assign fifo_intf_188.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_188;
    csv_file_dump cstatus_csv_dumper_188;
    df_fifo_monitor fifo_monitor_188;
    df_fifo_intf fifo_intf_189(clock,reset);
    assign fifo_intf_189.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_8_U.if_empty_n;
    assign fifo_intf_189.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_8_U.if_full_n;
    assign fifo_intf_189.fifo_rd_block = 0;
    assign fifo_intf_189.fifo_wr_block = 0;
    assign fifo_intf_189.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_189;
    csv_file_dump cstatus_csv_dumper_189;
    df_fifo_monitor fifo_monitor_189;
    df_fifo_intf fifo_intf_190(clock,reset);
    assign fifo_intf_190.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_8_U.if_empty_n;
    assign fifo_intf_190.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_8_U.if_full_n;
    assign fifo_intf_190.fifo_rd_block = 0;
    assign fifo_intf_190.fifo_wr_block = 0;
    assign fifo_intf_190.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_190;
    csv_file_dump cstatus_csv_dumper_190;
    df_fifo_monitor fifo_monitor_190;
    df_fifo_intf fifo_intf_191(clock,reset);
    assign fifo_intf_191.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_8_U.if_empty_n;
    assign fifo_intf_191.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_8_U.if_full_n;
    assign fifo_intf_191.fifo_rd_block = 0;
    assign fifo_intf_191.fifo_wr_block = 0;
    assign fifo_intf_191.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_191;
    csv_file_dump cstatus_csv_dumper_191;
    df_fifo_monitor fifo_monitor_191;
    df_fifo_intf fifo_intf_192(clock,reset);
    assign fifo_intf_192.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_8_U.if_empty_n;
    assign fifo_intf_192.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_8_U.if_full_n;
    assign fifo_intf_192.fifo_rd_block = 0;
    assign fifo_intf_192.fifo_wr_block = 0;
    assign fifo_intf_192.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_192;
    csv_file_dump cstatus_csv_dumper_192;
    df_fifo_monitor fifo_monitor_192;
    df_fifo_intf fifo_intf_193(clock,reset);
    assign fifo_intf_193.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_8_U.if_empty_n;
    assign fifo_intf_193.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_8_U.if_full_n;
    assign fifo_intf_193.fifo_rd_block = 0;
    assign fifo_intf_193.fifo_wr_block = 0;
    assign fifo_intf_193.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_193;
    csv_file_dump cstatus_csv_dumper_193;
    df_fifo_monitor fifo_monitor_193;
    df_fifo_intf fifo_intf_194(clock,reset);
    assign fifo_intf_194.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_8_U.if_empty_n;
    assign fifo_intf_194.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_8_U.if_full_n;
    assign fifo_intf_194.fifo_rd_block = 0;
    assign fifo_intf_194.fifo_wr_block = 0;
    assign fifo_intf_194.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_194;
    csv_file_dump cstatus_csv_dumper_194;
    df_fifo_monitor fifo_monitor_194;
    df_fifo_intf fifo_intf_195(clock,reset);
    assign fifo_intf_195.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_8_U.if_empty_n;
    assign fifo_intf_195.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_8_U.if_full_n;
    assign fifo_intf_195.fifo_rd_block = 0;
    assign fifo_intf_195.fifo_wr_block = 0;
    assign fifo_intf_195.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_195;
    csv_file_dump cstatus_csv_dumper_195;
    df_fifo_monitor fifo_monitor_195;
    df_fifo_intf fifo_intf_196(clock,reset);
    assign fifo_intf_196.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_8_U.if_empty_n;
    assign fifo_intf_196.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_8_U.if_full_n;
    assign fifo_intf_196.fifo_rd_block = 0;
    assign fifo_intf_196.fifo_wr_block = 0;
    assign fifo_intf_196.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_196;
    csv_file_dump cstatus_csv_dumper_196;
    df_fifo_monitor fifo_monitor_196;
    df_fifo_intf fifo_intf_197(clock,reset);
    assign fifo_intf_197.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_8_U.if_empty_n;
    assign fifo_intf_197.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_8_U.if_full_n;
    assign fifo_intf_197.fifo_rd_block = 0;
    assign fifo_intf_197.fifo_wr_block = 0;
    assign fifo_intf_197.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_197;
    csv_file_dump cstatus_csv_dumper_197;
    df_fifo_monitor fifo_monitor_197;
    df_fifo_intf fifo_intf_198(clock,reset);
    assign fifo_intf_198.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_8_U.if_empty_n;
    assign fifo_intf_198.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_8_U.if_full_n;
    assign fifo_intf_198.fifo_rd_block = 0;
    assign fifo_intf_198.fifo_wr_block = 0;
    assign fifo_intf_198.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_198;
    csv_file_dump cstatus_csv_dumper_198;
    df_fifo_monitor fifo_monitor_198;
    df_fifo_intf fifo_intf_199(clock,reset);
    assign fifo_intf_199.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_8_U.if_empty_n;
    assign fifo_intf_199.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_8_U.if_full_n;
    assign fifo_intf_199.fifo_rd_block = 0;
    assign fifo_intf_199.fifo_wr_block = 0;
    assign fifo_intf_199.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_199;
    csv_file_dump cstatus_csv_dumper_199;
    df_fifo_monitor fifo_monitor_199;
    df_fifo_intf fifo_intf_200(clock,reset);
    assign fifo_intf_200.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_8_U.if_empty_n;
    assign fifo_intf_200.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_8_U.if_full_n;
    assign fifo_intf_200.fifo_rd_block = 0;
    assign fifo_intf_200.fifo_wr_block = 0;
    assign fifo_intf_200.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_200;
    csv_file_dump cstatus_csv_dumper_200;
    df_fifo_monitor fifo_monitor_200;
    df_fifo_intf fifo_intf_201(clock,reset);
    assign fifo_intf_201.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_8_U.if_empty_n;
    assign fifo_intf_201.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_8_U.if_full_n;
    assign fifo_intf_201.fifo_rd_block = 0;
    assign fifo_intf_201.fifo_wr_block = 0;
    assign fifo_intf_201.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_201;
    csv_file_dump cstatus_csv_dumper_201;
    df_fifo_monitor fifo_monitor_201;
    df_fifo_intf fifo_intf_202(clock,reset);
    assign fifo_intf_202.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_8_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_8_U.if_empty_n;
    assign fifo_intf_202.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_8_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_8_U.if_full_n;
    assign fifo_intf_202.fifo_rd_block = 0;
    assign fifo_intf_202.fifo_wr_block = 0;
    assign fifo_intf_202.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_202;
    csv_file_dump cstatus_csv_dumper_202;
    df_fifo_monitor fifo_monitor_202;
    df_fifo_intf fifo_intf_203(clock,reset);
    assign fifo_intf_203.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_9_U.if_empty_n;
    assign fifo_intf_203.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_9_U.if_full_n;
    assign fifo_intf_203.fifo_rd_block = 0;
    assign fifo_intf_203.fifo_wr_block = 0;
    assign fifo_intf_203.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_203;
    csv_file_dump cstatus_csv_dumper_203;
    df_fifo_monitor fifo_monitor_203;
    df_fifo_intf fifo_intf_204(clock,reset);
    assign fifo_intf_204.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_9_U.if_empty_n;
    assign fifo_intf_204.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_9_U.if_full_n;
    assign fifo_intf_204.fifo_rd_block = 0;
    assign fifo_intf_204.fifo_wr_block = 0;
    assign fifo_intf_204.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_204;
    csv_file_dump cstatus_csv_dumper_204;
    df_fifo_monitor fifo_monitor_204;
    df_fifo_intf fifo_intf_205(clock,reset);
    assign fifo_intf_205.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_9_U.if_empty_n;
    assign fifo_intf_205.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_9_U.if_full_n;
    assign fifo_intf_205.fifo_rd_block = 0;
    assign fifo_intf_205.fifo_wr_block = 0;
    assign fifo_intf_205.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_205;
    csv_file_dump cstatus_csv_dumper_205;
    df_fifo_monitor fifo_monitor_205;
    df_fifo_intf fifo_intf_206(clock,reset);
    assign fifo_intf_206.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_9_U.if_empty_n;
    assign fifo_intf_206.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_9_U.if_full_n;
    assign fifo_intf_206.fifo_rd_block = 0;
    assign fifo_intf_206.fifo_wr_block = 0;
    assign fifo_intf_206.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_206;
    csv_file_dump cstatus_csv_dumper_206;
    df_fifo_monitor fifo_monitor_206;
    df_fifo_intf fifo_intf_207(clock,reset);
    assign fifo_intf_207.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_9_U.if_empty_n;
    assign fifo_intf_207.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_9_U.if_full_n;
    assign fifo_intf_207.fifo_rd_block = 0;
    assign fifo_intf_207.fifo_wr_block = 0;
    assign fifo_intf_207.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_207;
    csv_file_dump cstatus_csv_dumper_207;
    df_fifo_monitor fifo_monitor_207;
    df_fifo_intf fifo_intf_208(clock,reset);
    assign fifo_intf_208.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_9_U.if_empty_n;
    assign fifo_intf_208.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_9_U.if_full_n;
    assign fifo_intf_208.fifo_rd_block = 0;
    assign fifo_intf_208.fifo_wr_block = 0;
    assign fifo_intf_208.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_208;
    csv_file_dump cstatus_csv_dumper_208;
    df_fifo_monitor fifo_monitor_208;
    df_fifo_intf fifo_intf_209(clock,reset);
    assign fifo_intf_209.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_9_U.if_empty_n;
    assign fifo_intf_209.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_9_U.if_full_n;
    assign fifo_intf_209.fifo_rd_block = 0;
    assign fifo_intf_209.fifo_wr_block = 0;
    assign fifo_intf_209.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_209;
    csv_file_dump cstatus_csv_dumper_209;
    df_fifo_monitor fifo_monitor_209;
    df_fifo_intf fifo_intf_210(clock,reset);
    assign fifo_intf_210.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_9_U.if_empty_n;
    assign fifo_intf_210.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_9_U.if_full_n;
    assign fifo_intf_210.fifo_rd_block = 0;
    assign fifo_intf_210.fifo_wr_block = 0;
    assign fifo_intf_210.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_210;
    csv_file_dump cstatus_csv_dumper_210;
    df_fifo_monitor fifo_monitor_210;
    df_fifo_intf fifo_intf_211(clock,reset);
    assign fifo_intf_211.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_9_U.if_empty_n;
    assign fifo_intf_211.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_9_U.if_full_n;
    assign fifo_intf_211.fifo_rd_block = 0;
    assign fifo_intf_211.fifo_wr_block = 0;
    assign fifo_intf_211.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_211;
    csv_file_dump cstatus_csv_dumper_211;
    df_fifo_monitor fifo_monitor_211;
    df_fifo_intf fifo_intf_212(clock,reset);
    assign fifo_intf_212.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_9_U.if_empty_n;
    assign fifo_intf_212.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_9_U.if_full_n;
    assign fifo_intf_212.fifo_rd_block = 0;
    assign fifo_intf_212.fifo_wr_block = 0;
    assign fifo_intf_212.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_212;
    csv_file_dump cstatus_csv_dumper_212;
    df_fifo_monitor fifo_monitor_212;
    df_fifo_intf fifo_intf_213(clock,reset);
    assign fifo_intf_213.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_9_U.if_empty_n;
    assign fifo_intf_213.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_9_U.if_full_n;
    assign fifo_intf_213.fifo_rd_block = 0;
    assign fifo_intf_213.fifo_wr_block = 0;
    assign fifo_intf_213.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_213;
    csv_file_dump cstatus_csv_dumper_213;
    df_fifo_monitor fifo_monitor_213;
    df_fifo_intf fifo_intf_214(clock,reset);
    assign fifo_intf_214.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_9_U.if_empty_n;
    assign fifo_intf_214.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_9_U.if_full_n;
    assign fifo_intf_214.fifo_rd_block = 0;
    assign fifo_intf_214.fifo_wr_block = 0;
    assign fifo_intf_214.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_214;
    csv_file_dump cstatus_csv_dumper_214;
    df_fifo_monitor fifo_monitor_214;
    df_fifo_intf fifo_intf_215(clock,reset);
    assign fifo_intf_215.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_9_U.if_empty_n;
    assign fifo_intf_215.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_9_U.if_full_n;
    assign fifo_intf_215.fifo_rd_block = 0;
    assign fifo_intf_215.fifo_wr_block = 0;
    assign fifo_intf_215.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_215;
    csv_file_dump cstatus_csv_dumper_215;
    df_fifo_monitor fifo_monitor_215;
    df_fifo_intf fifo_intf_216(clock,reset);
    assign fifo_intf_216.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_9_U.if_empty_n;
    assign fifo_intf_216.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_9_U.if_full_n;
    assign fifo_intf_216.fifo_rd_block = 0;
    assign fifo_intf_216.fifo_wr_block = 0;
    assign fifo_intf_216.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_216;
    csv_file_dump cstatus_csv_dumper_216;
    df_fifo_monitor fifo_monitor_216;
    df_fifo_intf fifo_intf_217(clock,reset);
    assign fifo_intf_217.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_9_U.if_empty_n;
    assign fifo_intf_217.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_9_U.if_full_n;
    assign fifo_intf_217.fifo_rd_block = 0;
    assign fifo_intf_217.fifo_wr_block = 0;
    assign fifo_intf_217.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_217;
    csv_file_dump cstatus_csv_dumper_217;
    df_fifo_monitor fifo_monitor_217;
    df_fifo_intf fifo_intf_218(clock,reset);
    assign fifo_intf_218.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_9_U.if_empty_n;
    assign fifo_intf_218.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_9_U.if_full_n;
    assign fifo_intf_218.fifo_rd_block = 0;
    assign fifo_intf_218.fifo_wr_block = 0;
    assign fifo_intf_218.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_218;
    csv_file_dump cstatus_csv_dumper_218;
    df_fifo_monitor fifo_monitor_218;
    df_fifo_intf fifo_intf_219(clock,reset);
    assign fifo_intf_219.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_9_U.if_empty_n;
    assign fifo_intf_219.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_9_U.if_full_n;
    assign fifo_intf_219.fifo_rd_block = 0;
    assign fifo_intf_219.fifo_wr_block = 0;
    assign fifo_intf_219.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_219;
    csv_file_dump cstatus_csv_dumper_219;
    df_fifo_monitor fifo_monitor_219;
    df_fifo_intf fifo_intf_220(clock,reset);
    assign fifo_intf_220.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_9_U.if_empty_n;
    assign fifo_intf_220.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_9_U.if_full_n;
    assign fifo_intf_220.fifo_rd_block = 0;
    assign fifo_intf_220.fifo_wr_block = 0;
    assign fifo_intf_220.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_220;
    csv_file_dump cstatus_csv_dumper_220;
    df_fifo_monitor fifo_monitor_220;
    df_fifo_intf fifo_intf_221(clock,reset);
    assign fifo_intf_221.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_9_U.if_empty_n;
    assign fifo_intf_221.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_9_U.if_full_n;
    assign fifo_intf_221.fifo_rd_block = 0;
    assign fifo_intf_221.fifo_wr_block = 0;
    assign fifo_intf_221.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_221;
    csv_file_dump cstatus_csv_dumper_221;
    df_fifo_monitor fifo_monitor_221;
    df_fifo_intf fifo_intf_222(clock,reset);
    assign fifo_intf_222.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_9_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_9_U.if_empty_n;
    assign fifo_intf_222.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_9_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_9_U.if_full_n;
    assign fifo_intf_222.fifo_rd_block = 0;
    assign fifo_intf_222.fifo_wr_block = 0;
    assign fifo_intf_222.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_222;
    csv_file_dump cstatus_csv_dumper_222;
    df_fifo_monitor fifo_monitor_222;
    df_fifo_intf fifo_intf_223(clock,reset);
    assign fifo_intf_223.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_10_U.if_empty_n;
    assign fifo_intf_223.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_10_U.if_full_n;
    assign fifo_intf_223.fifo_rd_block = 0;
    assign fifo_intf_223.fifo_wr_block = 0;
    assign fifo_intf_223.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_223;
    csv_file_dump cstatus_csv_dumper_223;
    df_fifo_monitor fifo_monitor_223;
    df_fifo_intf fifo_intf_224(clock,reset);
    assign fifo_intf_224.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_10_U.if_empty_n;
    assign fifo_intf_224.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_10_U.if_full_n;
    assign fifo_intf_224.fifo_rd_block = 0;
    assign fifo_intf_224.fifo_wr_block = 0;
    assign fifo_intf_224.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_224;
    csv_file_dump cstatus_csv_dumper_224;
    df_fifo_monitor fifo_monitor_224;
    df_fifo_intf fifo_intf_225(clock,reset);
    assign fifo_intf_225.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_10_U.if_empty_n;
    assign fifo_intf_225.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_10_U.if_full_n;
    assign fifo_intf_225.fifo_rd_block = 0;
    assign fifo_intf_225.fifo_wr_block = 0;
    assign fifo_intf_225.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_225;
    csv_file_dump cstatus_csv_dumper_225;
    df_fifo_monitor fifo_monitor_225;
    df_fifo_intf fifo_intf_226(clock,reset);
    assign fifo_intf_226.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_10_U.if_empty_n;
    assign fifo_intf_226.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_10_U.if_full_n;
    assign fifo_intf_226.fifo_rd_block = 0;
    assign fifo_intf_226.fifo_wr_block = 0;
    assign fifo_intf_226.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_226;
    csv_file_dump cstatus_csv_dumper_226;
    df_fifo_monitor fifo_monitor_226;
    df_fifo_intf fifo_intf_227(clock,reset);
    assign fifo_intf_227.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_10_U.if_empty_n;
    assign fifo_intf_227.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_10_U.if_full_n;
    assign fifo_intf_227.fifo_rd_block = 0;
    assign fifo_intf_227.fifo_wr_block = 0;
    assign fifo_intf_227.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_227;
    csv_file_dump cstatus_csv_dumper_227;
    df_fifo_monitor fifo_monitor_227;
    df_fifo_intf fifo_intf_228(clock,reset);
    assign fifo_intf_228.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_10_U.if_empty_n;
    assign fifo_intf_228.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_10_U.if_full_n;
    assign fifo_intf_228.fifo_rd_block = 0;
    assign fifo_intf_228.fifo_wr_block = 0;
    assign fifo_intf_228.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_228;
    csv_file_dump cstatus_csv_dumper_228;
    df_fifo_monitor fifo_monitor_228;
    df_fifo_intf fifo_intf_229(clock,reset);
    assign fifo_intf_229.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_10_U.if_empty_n;
    assign fifo_intf_229.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_10_U.if_full_n;
    assign fifo_intf_229.fifo_rd_block = 0;
    assign fifo_intf_229.fifo_wr_block = 0;
    assign fifo_intf_229.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_229;
    csv_file_dump cstatus_csv_dumper_229;
    df_fifo_monitor fifo_monitor_229;
    df_fifo_intf fifo_intf_230(clock,reset);
    assign fifo_intf_230.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_10_U.if_empty_n;
    assign fifo_intf_230.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_10_U.if_full_n;
    assign fifo_intf_230.fifo_rd_block = 0;
    assign fifo_intf_230.fifo_wr_block = 0;
    assign fifo_intf_230.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_230;
    csv_file_dump cstatus_csv_dumper_230;
    df_fifo_monitor fifo_monitor_230;
    df_fifo_intf fifo_intf_231(clock,reset);
    assign fifo_intf_231.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_10_U.if_empty_n;
    assign fifo_intf_231.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_10_U.if_full_n;
    assign fifo_intf_231.fifo_rd_block = 0;
    assign fifo_intf_231.fifo_wr_block = 0;
    assign fifo_intf_231.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_231;
    csv_file_dump cstatus_csv_dumper_231;
    df_fifo_monitor fifo_monitor_231;
    df_fifo_intf fifo_intf_232(clock,reset);
    assign fifo_intf_232.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_10_U.if_empty_n;
    assign fifo_intf_232.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_10_U.if_full_n;
    assign fifo_intf_232.fifo_rd_block = 0;
    assign fifo_intf_232.fifo_wr_block = 0;
    assign fifo_intf_232.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_232;
    csv_file_dump cstatus_csv_dumper_232;
    df_fifo_monitor fifo_monitor_232;
    df_fifo_intf fifo_intf_233(clock,reset);
    assign fifo_intf_233.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_10_U.if_empty_n;
    assign fifo_intf_233.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_10_U.if_full_n;
    assign fifo_intf_233.fifo_rd_block = 0;
    assign fifo_intf_233.fifo_wr_block = 0;
    assign fifo_intf_233.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_233;
    csv_file_dump cstatus_csv_dumper_233;
    df_fifo_monitor fifo_monitor_233;
    df_fifo_intf fifo_intf_234(clock,reset);
    assign fifo_intf_234.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_10_U.if_empty_n;
    assign fifo_intf_234.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_10_U.if_full_n;
    assign fifo_intf_234.fifo_rd_block = 0;
    assign fifo_intf_234.fifo_wr_block = 0;
    assign fifo_intf_234.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_234;
    csv_file_dump cstatus_csv_dumper_234;
    df_fifo_monitor fifo_monitor_234;
    df_fifo_intf fifo_intf_235(clock,reset);
    assign fifo_intf_235.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_10_U.if_empty_n;
    assign fifo_intf_235.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_10_U.if_full_n;
    assign fifo_intf_235.fifo_rd_block = 0;
    assign fifo_intf_235.fifo_wr_block = 0;
    assign fifo_intf_235.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_235;
    csv_file_dump cstatus_csv_dumper_235;
    df_fifo_monitor fifo_monitor_235;
    df_fifo_intf fifo_intf_236(clock,reset);
    assign fifo_intf_236.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_10_U.if_empty_n;
    assign fifo_intf_236.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_10_U.if_full_n;
    assign fifo_intf_236.fifo_rd_block = 0;
    assign fifo_intf_236.fifo_wr_block = 0;
    assign fifo_intf_236.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_236;
    csv_file_dump cstatus_csv_dumper_236;
    df_fifo_monitor fifo_monitor_236;
    df_fifo_intf fifo_intf_237(clock,reset);
    assign fifo_intf_237.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_10_U.if_empty_n;
    assign fifo_intf_237.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_10_U.if_full_n;
    assign fifo_intf_237.fifo_rd_block = 0;
    assign fifo_intf_237.fifo_wr_block = 0;
    assign fifo_intf_237.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_237;
    csv_file_dump cstatus_csv_dumper_237;
    df_fifo_monitor fifo_monitor_237;
    df_fifo_intf fifo_intf_238(clock,reset);
    assign fifo_intf_238.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_10_U.if_empty_n;
    assign fifo_intf_238.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_10_U.if_full_n;
    assign fifo_intf_238.fifo_rd_block = 0;
    assign fifo_intf_238.fifo_wr_block = 0;
    assign fifo_intf_238.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_238;
    csv_file_dump cstatus_csv_dumper_238;
    df_fifo_monitor fifo_monitor_238;
    df_fifo_intf fifo_intf_239(clock,reset);
    assign fifo_intf_239.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_10_U.if_empty_n;
    assign fifo_intf_239.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_10_U.if_full_n;
    assign fifo_intf_239.fifo_rd_block = 0;
    assign fifo_intf_239.fifo_wr_block = 0;
    assign fifo_intf_239.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_239;
    csv_file_dump cstatus_csv_dumper_239;
    df_fifo_monitor fifo_monitor_239;
    df_fifo_intf fifo_intf_240(clock,reset);
    assign fifo_intf_240.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_10_U.if_empty_n;
    assign fifo_intf_240.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_10_U.if_full_n;
    assign fifo_intf_240.fifo_rd_block = 0;
    assign fifo_intf_240.fifo_wr_block = 0;
    assign fifo_intf_240.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_240;
    csv_file_dump cstatus_csv_dumper_240;
    df_fifo_monitor fifo_monitor_240;
    df_fifo_intf fifo_intf_241(clock,reset);
    assign fifo_intf_241.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_10_U.if_empty_n;
    assign fifo_intf_241.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_10_U.if_full_n;
    assign fifo_intf_241.fifo_rd_block = 0;
    assign fifo_intf_241.fifo_wr_block = 0;
    assign fifo_intf_241.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_241;
    csv_file_dump cstatus_csv_dumper_241;
    df_fifo_monitor fifo_monitor_241;
    df_fifo_intf fifo_intf_242(clock,reset);
    assign fifo_intf_242.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_10_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_10_U.if_empty_n;
    assign fifo_intf_242.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_10_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_10_U.if_full_n;
    assign fifo_intf_242.fifo_rd_block = 0;
    assign fifo_intf_242.fifo_wr_block = 0;
    assign fifo_intf_242.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_242;
    csv_file_dump cstatus_csv_dumper_242;
    df_fifo_monitor fifo_monitor_242;
    df_fifo_intf fifo_intf_243(clock,reset);
    assign fifo_intf_243.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_11_U.if_empty_n;
    assign fifo_intf_243.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_11_U.if_full_n;
    assign fifo_intf_243.fifo_rd_block = 0;
    assign fifo_intf_243.fifo_wr_block = 0;
    assign fifo_intf_243.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_243;
    csv_file_dump cstatus_csv_dumper_243;
    df_fifo_monitor fifo_monitor_243;
    df_fifo_intf fifo_intf_244(clock,reset);
    assign fifo_intf_244.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_11_U.if_empty_n;
    assign fifo_intf_244.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_11_U.if_full_n;
    assign fifo_intf_244.fifo_rd_block = 0;
    assign fifo_intf_244.fifo_wr_block = 0;
    assign fifo_intf_244.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_244;
    csv_file_dump cstatus_csv_dumper_244;
    df_fifo_monitor fifo_monitor_244;
    df_fifo_intf fifo_intf_245(clock,reset);
    assign fifo_intf_245.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_11_U.if_empty_n;
    assign fifo_intf_245.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_11_U.if_full_n;
    assign fifo_intf_245.fifo_rd_block = 0;
    assign fifo_intf_245.fifo_wr_block = 0;
    assign fifo_intf_245.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_245;
    csv_file_dump cstatus_csv_dumper_245;
    df_fifo_monitor fifo_monitor_245;
    df_fifo_intf fifo_intf_246(clock,reset);
    assign fifo_intf_246.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_11_U.if_empty_n;
    assign fifo_intf_246.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_11_U.if_full_n;
    assign fifo_intf_246.fifo_rd_block = 0;
    assign fifo_intf_246.fifo_wr_block = 0;
    assign fifo_intf_246.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_246;
    csv_file_dump cstatus_csv_dumper_246;
    df_fifo_monitor fifo_monitor_246;
    df_fifo_intf fifo_intf_247(clock,reset);
    assign fifo_intf_247.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_11_U.if_empty_n;
    assign fifo_intf_247.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_11_U.if_full_n;
    assign fifo_intf_247.fifo_rd_block = 0;
    assign fifo_intf_247.fifo_wr_block = 0;
    assign fifo_intf_247.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_247;
    csv_file_dump cstatus_csv_dumper_247;
    df_fifo_monitor fifo_monitor_247;
    df_fifo_intf fifo_intf_248(clock,reset);
    assign fifo_intf_248.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_11_U.if_empty_n;
    assign fifo_intf_248.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_11_U.if_full_n;
    assign fifo_intf_248.fifo_rd_block = 0;
    assign fifo_intf_248.fifo_wr_block = 0;
    assign fifo_intf_248.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_248;
    csv_file_dump cstatus_csv_dumper_248;
    df_fifo_monitor fifo_monitor_248;
    df_fifo_intf fifo_intf_249(clock,reset);
    assign fifo_intf_249.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_11_U.if_empty_n;
    assign fifo_intf_249.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_11_U.if_full_n;
    assign fifo_intf_249.fifo_rd_block = 0;
    assign fifo_intf_249.fifo_wr_block = 0;
    assign fifo_intf_249.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_249;
    csv_file_dump cstatus_csv_dumper_249;
    df_fifo_monitor fifo_monitor_249;
    df_fifo_intf fifo_intf_250(clock,reset);
    assign fifo_intf_250.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_11_U.if_empty_n;
    assign fifo_intf_250.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_11_U.if_full_n;
    assign fifo_intf_250.fifo_rd_block = 0;
    assign fifo_intf_250.fifo_wr_block = 0;
    assign fifo_intf_250.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_250;
    csv_file_dump cstatus_csv_dumper_250;
    df_fifo_monitor fifo_monitor_250;
    df_fifo_intf fifo_intf_251(clock,reset);
    assign fifo_intf_251.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_11_U.if_empty_n;
    assign fifo_intf_251.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_11_U.if_full_n;
    assign fifo_intf_251.fifo_rd_block = 0;
    assign fifo_intf_251.fifo_wr_block = 0;
    assign fifo_intf_251.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_251;
    csv_file_dump cstatus_csv_dumper_251;
    df_fifo_monitor fifo_monitor_251;
    df_fifo_intf fifo_intf_252(clock,reset);
    assign fifo_intf_252.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_11_U.if_empty_n;
    assign fifo_intf_252.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_11_U.if_full_n;
    assign fifo_intf_252.fifo_rd_block = 0;
    assign fifo_intf_252.fifo_wr_block = 0;
    assign fifo_intf_252.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_252;
    csv_file_dump cstatus_csv_dumper_252;
    df_fifo_monitor fifo_monitor_252;
    df_fifo_intf fifo_intf_253(clock,reset);
    assign fifo_intf_253.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_11_U.if_empty_n;
    assign fifo_intf_253.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_11_U.if_full_n;
    assign fifo_intf_253.fifo_rd_block = 0;
    assign fifo_intf_253.fifo_wr_block = 0;
    assign fifo_intf_253.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_253;
    csv_file_dump cstatus_csv_dumper_253;
    df_fifo_monitor fifo_monitor_253;
    df_fifo_intf fifo_intf_254(clock,reset);
    assign fifo_intf_254.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_11_U.if_empty_n;
    assign fifo_intf_254.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_11_U.if_full_n;
    assign fifo_intf_254.fifo_rd_block = 0;
    assign fifo_intf_254.fifo_wr_block = 0;
    assign fifo_intf_254.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_254;
    csv_file_dump cstatus_csv_dumper_254;
    df_fifo_monitor fifo_monitor_254;
    df_fifo_intf fifo_intf_255(clock,reset);
    assign fifo_intf_255.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_11_U.if_empty_n;
    assign fifo_intf_255.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_11_U.if_full_n;
    assign fifo_intf_255.fifo_rd_block = 0;
    assign fifo_intf_255.fifo_wr_block = 0;
    assign fifo_intf_255.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_255;
    csv_file_dump cstatus_csv_dumper_255;
    df_fifo_monitor fifo_monitor_255;
    df_fifo_intf fifo_intf_256(clock,reset);
    assign fifo_intf_256.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_11_U.if_empty_n;
    assign fifo_intf_256.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_11_U.if_full_n;
    assign fifo_intf_256.fifo_rd_block = 0;
    assign fifo_intf_256.fifo_wr_block = 0;
    assign fifo_intf_256.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_256;
    csv_file_dump cstatus_csv_dumper_256;
    df_fifo_monitor fifo_monitor_256;
    df_fifo_intf fifo_intf_257(clock,reset);
    assign fifo_intf_257.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_11_U.if_empty_n;
    assign fifo_intf_257.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_11_U.if_full_n;
    assign fifo_intf_257.fifo_rd_block = 0;
    assign fifo_intf_257.fifo_wr_block = 0;
    assign fifo_intf_257.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_257;
    csv_file_dump cstatus_csv_dumper_257;
    df_fifo_monitor fifo_monitor_257;
    df_fifo_intf fifo_intf_258(clock,reset);
    assign fifo_intf_258.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_11_U.if_empty_n;
    assign fifo_intf_258.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_11_U.if_full_n;
    assign fifo_intf_258.fifo_rd_block = 0;
    assign fifo_intf_258.fifo_wr_block = 0;
    assign fifo_intf_258.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_258;
    csv_file_dump cstatus_csv_dumper_258;
    df_fifo_monitor fifo_monitor_258;
    df_fifo_intf fifo_intf_259(clock,reset);
    assign fifo_intf_259.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_11_U.if_empty_n;
    assign fifo_intf_259.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_11_U.if_full_n;
    assign fifo_intf_259.fifo_rd_block = 0;
    assign fifo_intf_259.fifo_wr_block = 0;
    assign fifo_intf_259.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_259;
    csv_file_dump cstatus_csv_dumper_259;
    df_fifo_monitor fifo_monitor_259;
    df_fifo_intf fifo_intf_260(clock,reset);
    assign fifo_intf_260.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_11_U.if_empty_n;
    assign fifo_intf_260.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_11_U.if_full_n;
    assign fifo_intf_260.fifo_rd_block = 0;
    assign fifo_intf_260.fifo_wr_block = 0;
    assign fifo_intf_260.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_260;
    csv_file_dump cstatus_csv_dumper_260;
    df_fifo_monitor fifo_monitor_260;
    df_fifo_intf fifo_intf_261(clock,reset);
    assign fifo_intf_261.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_11_U.if_empty_n;
    assign fifo_intf_261.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_11_U.if_full_n;
    assign fifo_intf_261.fifo_rd_block = 0;
    assign fifo_intf_261.fifo_wr_block = 0;
    assign fifo_intf_261.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_261;
    csv_file_dump cstatus_csv_dumper_261;
    df_fifo_monitor fifo_monitor_261;
    df_fifo_intf fifo_intf_262(clock,reset);
    assign fifo_intf_262.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_11_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_11_U.if_empty_n;
    assign fifo_intf_262.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_11_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_11_U.if_full_n;
    assign fifo_intf_262.fifo_rd_block = 0;
    assign fifo_intf_262.fifo_wr_block = 0;
    assign fifo_intf_262.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_262;
    csv_file_dump cstatus_csv_dumper_262;
    df_fifo_monitor fifo_monitor_262;
    df_fifo_intf fifo_intf_263(clock,reset);
    assign fifo_intf_263.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_12_U.if_empty_n;
    assign fifo_intf_263.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_12_U.if_full_n;
    assign fifo_intf_263.fifo_rd_block = 0;
    assign fifo_intf_263.fifo_wr_block = 0;
    assign fifo_intf_263.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_263;
    csv_file_dump cstatus_csv_dumper_263;
    df_fifo_monitor fifo_monitor_263;
    df_fifo_intf fifo_intf_264(clock,reset);
    assign fifo_intf_264.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_12_U.if_empty_n;
    assign fifo_intf_264.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_12_U.if_full_n;
    assign fifo_intf_264.fifo_rd_block = 0;
    assign fifo_intf_264.fifo_wr_block = 0;
    assign fifo_intf_264.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_264;
    csv_file_dump cstatus_csv_dumper_264;
    df_fifo_monitor fifo_monitor_264;
    df_fifo_intf fifo_intf_265(clock,reset);
    assign fifo_intf_265.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_12_U.if_empty_n;
    assign fifo_intf_265.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_12_U.if_full_n;
    assign fifo_intf_265.fifo_rd_block = 0;
    assign fifo_intf_265.fifo_wr_block = 0;
    assign fifo_intf_265.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_265;
    csv_file_dump cstatus_csv_dumper_265;
    df_fifo_monitor fifo_monitor_265;
    df_fifo_intf fifo_intf_266(clock,reset);
    assign fifo_intf_266.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_12_U.if_empty_n;
    assign fifo_intf_266.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_12_U.if_full_n;
    assign fifo_intf_266.fifo_rd_block = 0;
    assign fifo_intf_266.fifo_wr_block = 0;
    assign fifo_intf_266.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_266;
    csv_file_dump cstatus_csv_dumper_266;
    df_fifo_monitor fifo_monitor_266;
    df_fifo_intf fifo_intf_267(clock,reset);
    assign fifo_intf_267.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_12_U.if_empty_n;
    assign fifo_intf_267.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_12_U.if_full_n;
    assign fifo_intf_267.fifo_rd_block = 0;
    assign fifo_intf_267.fifo_wr_block = 0;
    assign fifo_intf_267.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_267;
    csv_file_dump cstatus_csv_dumper_267;
    df_fifo_monitor fifo_monitor_267;
    df_fifo_intf fifo_intf_268(clock,reset);
    assign fifo_intf_268.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_12_U.if_empty_n;
    assign fifo_intf_268.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_12_U.if_full_n;
    assign fifo_intf_268.fifo_rd_block = 0;
    assign fifo_intf_268.fifo_wr_block = 0;
    assign fifo_intf_268.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_268;
    csv_file_dump cstatus_csv_dumper_268;
    df_fifo_monitor fifo_monitor_268;
    df_fifo_intf fifo_intf_269(clock,reset);
    assign fifo_intf_269.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_12_U.if_empty_n;
    assign fifo_intf_269.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_12_U.if_full_n;
    assign fifo_intf_269.fifo_rd_block = 0;
    assign fifo_intf_269.fifo_wr_block = 0;
    assign fifo_intf_269.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_269;
    csv_file_dump cstatus_csv_dumper_269;
    df_fifo_monitor fifo_monitor_269;
    df_fifo_intf fifo_intf_270(clock,reset);
    assign fifo_intf_270.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_12_U.if_empty_n;
    assign fifo_intf_270.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_12_U.if_full_n;
    assign fifo_intf_270.fifo_rd_block = 0;
    assign fifo_intf_270.fifo_wr_block = 0;
    assign fifo_intf_270.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_270;
    csv_file_dump cstatus_csv_dumper_270;
    df_fifo_monitor fifo_monitor_270;
    df_fifo_intf fifo_intf_271(clock,reset);
    assign fifo_intf_271.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_12_U.if_empty_n;
    assign fifo_intf_271.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_12_U.if_full_n;
    assign fifo_intf_271.fifo_rd_block = 0;
    assign fifo_intf_271.fifo_wr_block = 0;
    assign fifo_intf_271.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_271;
    csv_file_dump cstatus_csv_dumper_271;
    df_fifo_monitor fifo_monitor_271;
    df_fifo_intf fifo_intf_272(clock,reset);
    assign fifo_intf_272.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_12_U.if_empty_n;
    assign fifo_intf_272.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_12_U.if_full_n;
    assign fifo_intf_272.fifo_rd_block = 0;
    assign fifo_intf_272.fifo_wr_block = 0;
    assign fifo_intf_272.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_272;
    csv_file_dump cstatus_csv_dumper_272;
    df_fifo_monitor fifo_monitor_272;
    df_fifo_intf fifo_intf_273(clock,reset);
    assign fifo_intf_273.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_12_U.if_empty_n;
    assign fifo_intf_273.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_12_U.if_full_n;
    assign fifo_intf_273.fifo_rd_block = 0;
    assign fifo_intf_273.fifo_wr_block = 0;
    assign fifo_intf_273.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_273;
    csv_file_dump cstatus_csv_dumper_273;
    df_fifo_monitor fifo_monitor_273;
    df_fifo_intf fifo_intf_274(clock,reset);
    assign fifo_intf_274.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_12_U.if_empty_n;
    assign fifo_intf_274.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_12_U.if_full_n;
    assign fifo_intf_274.fifo_rd_block = 0;
    assign fifo_intf_274.fifo_wr_block = 0;
    assign fifo_intf_274.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_274;
    csv_file_dump cstatus_csv_dumper_274;
    df_fifo_monitor fifo_monitor_274;
    df_fifo_intf fifo_intf_275(clock,reset);
    assign fifo_intf_275.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_12_U.if_empty_n;
    assign fifo_intf_275.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_12_U.if_full_n;
    assign fifo_intf_275.fifo_rd_block = 0;
    assign fifo_intf_275.fifo_wr_block = 0;
    assign fifo_intf_275.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_275;
    csv_file_dump cstatus_csv_dumper_275;
    df_fifo_monitor fifo_monitor_275;
    df_fifo_intf fifo_intf_276(clock,reset);
    assign fifo_intf_276.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_12_U.if_empty_n;
    assign fifo_intf_276.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_12_U.if_full_n;
    assign fifo_intf_276.fifo_rd_block = 0;
    assign fifo_intf_276.fifo_wr_block = 0;
    assign fifo_intf_276.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_276;
    csv_file_dump cstatus_csv_dumper_276;
    df_fifo_monitor fifo_monitor_276;
    df_fifo_intf fifo_intf_277(clock,reset);
    assign fifo_intf_277.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_12_U.if_empty_n;
    assign fifo_intf_277.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_12_U.if_full_n;
    assign fifo_intf_277.fifo_rd_block = 0;
    assign fifo_intf_277.fifo_wr_block = 0;
    assign fifo_intf_277.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_277;
    csv_file_dump cstatus_csv_dumper_277;
    df_fifo_monitor fifo_monitor_277;
    df_fifo_intf fifo_intf_278(clock,reset);
    assign fifo_intf_278.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_12_U.if_empty_n;
    assign fifo_intf_278.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_12_U.if_full_n;
    assign fifo_intf_278.fifo_rd_block = 0;
    assign fifo_intf_278.fifo_wr_block = 0;
    assign fifo_intf_278.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_278;
    csv_file_dump cstatus_csv_dumper_278;
    df_fifo_monitor fifo_monitor_278;
    df_fifo_intf fifo_intf_279(clock,reset);
    assign fifo_intf_279.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_12_U.if_empty_n;
    assign fifo_intf_279.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_12_U.if_full_n;
    assign fifo_intf_279.fifo_rd_block = 0;
    assign fifo_intf_279.fifo_wr_block = 0;
    assign fifo_intf_279.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_279;
    csv_file_dump cstatus_csv_dumper_279;
    df_fifo_monitor fifo_monitor_279;
    df_fifo_intf fifo_intf_280(clock,reset);
    assign fifo_intf_280.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_12_U.if_empty_n;
    assign fifo_intf_280.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_12_U.if_full_n;
    assign fifo_intf_280.fifo_rd_block = 0;
    assign fifo_intf_280.fifo_wr_block = 0;
    assign fifo_intf_280.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_280;
    csv_file_dump cstatus_csv_dumper_280;
    df_fifo_monitor fifo_monitor_280;
    df_fifo_intf fifo_intf_281(clock,reset);
    assign fifo_intf_281.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_12_U.if_empty_n;
    assign fifo_intf_281.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_12_U.if_full_n;
    assign fifo_intf_281.fifo_rd_block = 0;
    assign fifo_intf_281.fifo_wr_block = 0;
    assign fifo_intf_281.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_281;
    csv_file_dump cstatus_csv_dumper_281;
    df_fifo_monitor fifo_monitor_281;
    df_fifo_intf fifo_intf_282(clock,reset);
    assign fifo_intf_282.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_12_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_12_U.if_empty_n;
    assign fifo_intf_282.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_12_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_12_U.if_full_n;
    assign fifo_intf_282.fifo_rd_block = 0;
    assign fifo_intf_282.fifo_wr_block = 0;
    assign fifo_intf_282.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_282;
    csv_file_dump cstatus_csv_dumper_282;
    df_fifo_monitor fifo_monitor_282;
    df_fifo_intf fifo_intf_283(clock,reset);
    assign fifo_intf_283.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_13_U.if_empty_n;
    assign fifo_intf_283.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_13_U.if_full_n;
    assign fifo_intf_283.fifo_rd_block = 0;
    assign fifo_intf_283.fifo_wr_block = 0;
    assign fifo_intf_283.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_283;
    csv_file_dump cstatus_csv_dumper_283;
    df_fifo_monitor fifo_monitor_283;
    df_fifo_intf fifo_intf_284(clock,reset);
    assign fifo_intf_284.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_13_U.if_empty_n;
    assign fifo_intf_284.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_13_U.if_full_n;
    assign fifo_intf_284.fifo_rd_block = 0;
    assign fifo_intf_284.fifo_wr_block = 0;
    assign fifo_intf_284.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_284;
    csv_file_dump cstatus_csv_dumper_284;
    df_fifo_monitor fifo_monitor_284;
    df_fifo_intf fifo_intf_285(clock,reset);
    assign fifo_intf_285.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_13_U.if_empty_n;
    assign fifo_intf_285.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_13_U.if_full_n;
    assign fifo_intf_285.fifo_rd_block = 0;
    assign fifo_intf_285.fifo_wr_block = 0;
    assign fifo_intf_285.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_285;
    csv_file_dump cstatus_csv_dumper_285;
    df_fifo_monitor fifo_monitor_285;
    df_fifo_intf fifo_intf_286(clock,reset);
    assign fifo_intf_286.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_13_U.if_empty_n;
    assign fifo_intf_286.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_13_U.if_full_n;
    assign fifo_intf_286.fifo_rd_block = 0;
    assign fifo_intf_286.fifo_wr_block = 0;
    assign fifo_intf_286.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_286;
    csv_file_dump cstatus_csv_dumper_286;
    df_fifo_monitor fifo_monitor_286;
    df_fifo_intf fifo_intf_287(clock,reset);
    assign fifo_intf_287.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_13_U.if_empty_n;
    assign fifo_intf_287.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_13_U.if_full_n;
    assign fifo_intf_287.fifo_rd_block = 0;
    assign fifo_intf_287.fifo_wr_block = 0;
    assign fifo_intf_287.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_287;
    csv_file_dump cstatus_csv_dumper_287;
    df_fifo_monitor fifo_monitor_287;
    df_fifo_intf fifo_intf_288(clock,reset);
    assign fifo_intf_288.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_13_U.if_empty_n;
    assign fifo_intf_288.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_13_U.if_full_n;
    assign fifo_intf_288.fifo_rd_block = 0;
    assign fifo_intf_288.fifo_wr_block = 0;
    assign fifo_intf_288.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_288;
    csv_file_dump cstatus_csv_dumper_288;
    df_fifo_monitor fifo_monitor_288;
    df_fifo_intf fifo_intf_289(clock,reset);
    assign fifo_intf_289.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_13_U.if_empty_n;
    assign fifo_intf_289.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_13_U.if_full_n;
    assign fifo_intf_289.fifo_rd_block = 0;
    assign fifo_intf_289.fifo_wr_block = 0;
    assign fifo_intf_289.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_289;
    csv_file_dump cstatus_csv_dumper_289;
    df_fifo_monitor fifo_monitor_289;
    df_fifo_intf fifo_intf_290(clock,reset);
    assign fifo_intf_290.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_13_U.if_empty_n;
    assign fifo_intf_290.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_13_U.if_full_n;
    assign fifo_intf_290.fifo_rd_block = 0;
    assign fifo_intf_290.fifo_wr_block = 0;
    assign fifo_intf_290.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_290;
    csv_file_dump cstatus_csv_dumper_290;
    df_fifo_monitor fifo_monitor_290;
    df_fifo_intf fifo_intf_291(clock,reset);
    assign fifo_intf_291.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_13_U.if_empty_n;
    assign fifo_intf_291.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_13_U.if_full_n;
    assign fifo_intf_291.fifo_rd_block = 0;
    assign fifo_intf_291.fifo_wr_block = 0;
    assign fifo_intf_291.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_291;
    csv_file_dump cstatus_csv_dumper_291;
    df_fifo_monitor fifo_monitor_291;
    df_fifo_intf fifo_intf_292(clock,reset);
    assign fifo_intf_292.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_13_U.if_empty_n;
    assign fifo_intf_292.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_13_U.if_full_n;
    assign fifo_intf_292.fifo_rd_block = 0;
    assign fifo_intf_292.fifo_wr_block = 0;
    assign fifo_intf_292.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_292;
    csv_file_dump cstatus_csv_dumper_292;
    df_fifo_monitor fifo_monitor_292;
    df_fifo_intf fifo_intf_293(clock,reset);
    assign fifo_intf_293.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_13_U.if_empty_n;
    assign fifo_intf_293.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_13_U.if_full_n;
    assign fifo_intf_293.fifo_rd_block = 0;
    assign fifo_intf_293.fifo_wr_block = 0;
    assign fifo_intf_293.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_293;
    csv_file_dump cstatus_csv_dumper_293;
    df_fifo_monitor fifo_monitor_293;
    df_fifo_intf fifo_intf_294(clock,reset);
    assign fifo_intf_294.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_13_U.if_empty_n;
    assign fifo_intf_294.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_13_U.if_full_n;
    assign fifo_intf_294.fifo_rd_block = 0;
    assign fifo_intf_294.fifo_wr_block = 0;
    assign fifo_intf_294.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_294;
    csv_file_dump cstatus_csv_dumper_294;
    df_fifo_monitor fifo_monitor_294;
    df_fifo_intf fifo_intf_295(clock,reset);
    assign fifo_intf_295.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_13_U.if_empty_n;
    assign fifo_intf_295.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_13_U.if_full_n;
    assign fifo_intf_295.fifo_rd_block = 0;
    assign fifo_intf_295.fifo_wr_block = 0;
    assign fifo_intf_295.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_295;
    csv_file_dump cstatus_csv_dumper_295;
    df_fifo_monitor fifo_monitor_295;
    df_fifo_intf fifo_intf_296(clock,reset);
    assign fifo_intf_296.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_13_U.if_empty_n;
    assign fifo_intf_296.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_13_U.if_full_n;
    assign fifo_intf_296.fifo_rd_block = 0;
    assign fifo_intf_296.fifo_wr_block = 0;
    assign fifo_intf_296.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_296;
    csv_file_dump cstatus_csv_dumper_296;
    df_fifo_monitor fifo_monitor_296;
    df_fifo_intf fifo_intf_297(clock,reset);
    assign fifo_intf_297.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_13_U.if_empty_n;
    assign fifo_intf_297.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_13_U.if_full_n;
    assign fifo_intf_297.fifo_rd_block = 0;
    assign fifo_intf_297.fifo_wr_block = 0;
    assign fifo_intf_297.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_297;
    csv_file_dump cstatus_csv_dumper_297;
    df_fifo_monitor fifo_monitor_297;
    df_fifo_intf fifo_intf_298(clock,reset);
    assign fifo_intf_298.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_13_U.if_empty_n;
    assign fifo_intf_298.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_13_U.if_full_n;
    assign fifo_intf_298.fifo_rd_block = 0;
    assign fifo_intf_298.fifo_wr_block = 0;
    assign fifo_intf_298.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_298;
    csv_file_dump cstatus_csv_dumper_298;
    df_fifo_monitor fifo_monitor_298;
    df_fifo_intf fifo_intf_299(clock,reset);
    assign fifo_intf_299.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_13_U.if_empty_n;
    assign fifo_intf_299.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_13_U.if_full_n;
    assign fifo_intf_299.fifo_rd_block = 0;
    assign fifo_intf_299.fifo_wr_block = 0;
    assign fifo_intf_299.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_299;
    csv_file_dump cstatus_csv_dumper_299;
    df_fifo_monitor fifo_monitor_299;
    df_fifo_intf fifo_intf_300(clock,reset);
    assign fifo_intf_300.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_13_U.if_empty_n;
    assign fifo_intf_300.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_13_U.if_full_n;
    assign fifo_intf_300.fifo_rd_block = 0;
    assign fifo_intf_300.fifo_wr_block = 0;
    assign fifo_intf_300.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_300;
    csv_file_dump cstatus_csv_dumper_300;
    df_fifo_monitor fifo_monitor_300;
    df_fifo_intf fifo_intf_301(clock,reset);
    assign fifo_intf_301.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_13_U.if_empty_n;
    assign fifo_intf_301.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_13_U.if_full_n;
    assign fifo_intf_301.fifo_rd_block = 0;
    assign fifo_intf_301.fifo_wr_block = 0;
    assign fifo_intf_301.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_301;
    csv_file_dump cstatus_csv_dumper_301;
    df_fifo_monitor fifo_monitor_301;
    df_fifo_intf fifo_intf_302(clock,reset);
    assign fifo_intf_302.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_13_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_13_U.if_empty_n;
    assign fifo_intf_302.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_13_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_13_U.if_full_n;
    assign fifo_intf_302.fifo_rd_block = 0;
    assign fifo_intf_302.fifo_wr_block = 0;
    assign fifo_intf_302.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_302;
    csv_file_dump cstatus_csv_dumper_302;
    df_fifo_monitor fifo_monitor_302;
    df_fifo_intf fifo_intf_303(clock,reset);
    assign fifo_intf_303.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_14_U.if_empty_n;
    assign fifo_intf_303.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_14_U.if_full_n;
    assign fifo_intf_303.fifo_rd_block = 0;
    assign fifo_intf_303.fifo_wr_block = 0;
    assign fifo_intf_303.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_303;
    csv_file_dump cstatus_csv_dumper_303;
    df_fifo_monitor fifo_monitor_303;
    df_fifo_intf fifo_intf_304(clock,reset);
    assign fifo_intf_304.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_14_U.if_empty_n;
    assign fifo_intf_304.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_14_U.if_full_n;
    assign fifo_intf_304.fifo_rd_block = 0;
    assign fifo_intf_304.fifo_wr_block = 0;
    assign fifo_intf_304.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_304;
    csv_file_dump cstatus_csv_dumper_304;
    df_fifo_monitor fifo_monitor_304;
    df_fifo_intf fifo_intf_305(clock,reset);
    assign fifo_intf_305.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_14_U.if_empty_n;
    assign fifo_intf_305.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_14_U.if_full_n;
    assign fifo_intf_305.fifo_rd_block = 0;
    assign fifo_intf_305.fifo_wr_block = 0;
    assign fifo_intf_305.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_305;
    csv_file_dump cstatus_csv_dumper_305;
    df_fifo_monitor fifo_monitor_305;
    df_fifo_intf fifo_intf_306(clock,reset);
    assign fifo_intf_306.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_14_U.if_empty_n;
    assign fifo_intf_306.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_14_U.if_full_n;
    assign fifo_intf_306.fifo_rd_block = 0;
    assign fifo_intf_306.fifo_wr_block = 0;
    assign fifo_intf_306.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_306;
    csv_file_dump cstatus_csv_dumper_306;
    df_fifo_monitor fifo_monitor_306;
    df_fifo_intf fifo_intf_307(clock,reset);
    assign fifo_intf_307.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_14_U.if_empty_n;
    assign fifo_intf_307.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_14_U.if_full_n;
    assign fifo_intf_307.fifo_rd_block = 0;
    assign fifo_intf_307.fifo_wr_block = 0;
    assign fifo_intf_307.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_307;
    csv_file_dump cstatus_csv_dumper_307;
    df_fifo_monitor fifo_monitor_307;
    df_fifo_intf fifo_intf_308(clock,reset);
    assign fifo_intf_308.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_14_U.if_empty_n;
    assign fifo_intf_308.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_14_U.if_full_n;
    assign fifo_intf_308.fifo_rd_block = 0;
    assign fifo_intf_308.fifo_wr_block = 0;
    assign fifo_intf_308.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_308;
    csv_file_dump cstatus_csv_dumper_308;
    df_fifo_monitor fifo_monitor_308;
    df_fifo_intf fifo_intf_309(clock,reset);
    assign fifo_intf_309.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_14_U.if_empty_n;
    assign fifo_intf_309.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_14_U.if_full_n;
    assign fifo_intf_309.fifo_rd_block = 0;
    assign fifo_intf_309.fifo_wr_block = 0;
    assign fifo_intf_309.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_309;
    csv_file_dump cstatus_csv_dumper_309;
    df_fifo_monitor fifo_monitor_309;
    df_fifo_intf fifo_intf_310(clock,reset);
    assign fifo_intf_310.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_14_U.if_empty_n;
    assign fifo_intf_310.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_14_U.if_full_n;
    assign fifo_intf_310.fifo_rd_block = 0;
    assign fifo_intf_310.fifo_wr_block = 0;
    assign fifo_intf_310.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_310;
    csv_file_dump cstatus_csv_dumper_310;
    df_fifo_monitor fifo_monitor_310;
    df_fifo_intf fifo_intf_311(clock,reset);
    assign fifo_intf_311.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_14_U.if_empty_n;
    assign fifo_intf_311.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_14_U.if_full_n;
    assign fifo_intf_311.fifo_rd_block = 0;
    assign fifo_intf_311.fifo_wr_block = 0;
    assign fifo_intf_311.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_311;
    csv_file_dump cstatus_csv_dumper_311;
    df_fifo_monitor fifo_monitor_311;
    df_fifo_intf fifo_intf_312(clock,reset);
    assign fifo_intf_312.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_14_U.if_empty_n;
    assign fifo_intf_312.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_14_U.if_full_n;
    assign fifo_intf_312.fifo_rd_block = 0;
    assign fifo_intf_312.fifo_wr_block = 0;
    assign fifo_intf_312.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_312;
    csv_file_dump cstatus_csv_dumper_312;
    df_fifo_monitor fifo_monitor_312;
    df_fifo_intf fifo_intf_313(clock,reset);
    assign fifo_intf_313.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_14_U.if_empty_n;
    assign fifo_intf_313.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_14_U.if_full_n;
    assign fifo_intf_313.fifo_rd_block = 0;
    assign fifo_intf_313.fifo_wr_block = 0;
    assign fifo_intf_313.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_313;
    csv_file_dump cstatus_csv_dumper_313;
    df_fifo_monitor fifo_monitor_313;
    df_fifo_intf fifo_intf_314(clock,reset);
    assign fifo_intf_314.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_14_U.if_empty_n;
    assign fifo_intf_314.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_14_U.if_full_n;
    assign fifo_intf_314.fifo_rd_block = 0;
    assign fifo_intf_314.fifo_wr_block = 0;
    assign fifo_intf_314.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_314;
    csv_file_dump cstatus_csv_dumper_314;
    df_fifo_monitor fifo_monitor_314;
    df_fifo_intf fifo_intf_315(clock,reset);
    assign fifo_intf_315.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_14_U.if_empty_n;
    assign fifo_intf_315.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_14_U.if_full_n;
    assign fifo_intf_315.fifo_rd_block = 0;
    assign fifo_intf_315.fifo_wr_block = 0;
    assign fifo_intf_315.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_315;
    csv_file_dump cstatus_csv_dumper_315;
    df_fifo_monitor fifo_monitor_315;
    df_fifo_intf fifo_intf_316(clock,reset);
    assign fifo_intf_316.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_14_U.if_empty_n;
    assign fifo_intf_316.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_14_U.if_full_n;
    assign fifo_intf_316.fifo_rd_block = 0;
    assign fifo_intf_316.fifo_wr_block = 0;
    assign fifo_intf_316.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_316;
    csv_file_dump cstatus_csv_dumper_316;
    df_fifo_monitor fifo_monitor_316;
    df_fifo_intf fifo_intf_317(clock,reset);
    assign fifo_intf_317.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_14_U.if_empty_n;
    assign fifo_intf_317.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_14_U.if_full_n;
    assign fifo_intf_317.fifo_rd_block = 0;
    assign fifo_intf_317.fifo_wr_block = 0;
    assign fifo_intf_317.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_317;
    csv_file_dump cstatus_csv_dumper_317;
    df_fifo_monitor fifo_monitor_317;
    df_fifo_intf fifo_intf_318(clock,reset);
    assign fifo_intf_318.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_14_U.if_empty_n;
    assign fifo_intf_318.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_14_U.if_full_n;
    assign fifo_intf_318.fifo_rd_block = 0;
    assign fifo_intf_318.fifo_wr_block = 0;
    assign fifo_intf_318.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_318;
    csv_file_dump cstatus_csv_dumper_318;
    df_fifo_monitor fifo_monitor_318;
    df_fifo_intf fifo_intf_319(clock,reset);
    assign fifo_intf_319.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_14_U.if_empty_n;
    assign fifo_intf_319.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_14_U.if_full_n;
    assign fifo_intf_319.fifo_rd_block = 0;
    assign fifo_intf_319.fifo_wr_block = 0;
    assign fifo_intf_319.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_319;
    csv_file_dump cstatus_csv_dumper_319;
    df_fifo_monitor fifo_monitor_319;
    df_fifo_intf fifo_intf_320(clock,reset);
    assign fifo_intf_320.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_14_U.if_empty_n;
    assign fifo_intf_320.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_14_U.if_full_n;
    assign fifo_intf_320.fifo_rd_block = 0;
    assign fifo_intf_320.fifo_wr_block = 0;
    assign fifo_intf_320.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_320;
    csv_file_dump cstatus_csv_dumper_320;
    df_fifo_monitor fifo_monitor_320;
    df_fifo_intf fifo_intf_321(clock,reset);
    assign fifo_intf_321.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_14_U.if_empty_n;
    assign fifo_intf_321.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_14_U.if_full_n;
    assign fifo_intf_321.fifo_rd_block = 0;
    assign fifo_intf_321.fifo_wr_block = 0;
    assign fifo_intf_321.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_321;
    csv_file_dump cstatus_csv_dumper_321;
    df_fifo_monitor fifo_monitor_321;
    df_fifo_intf fifo_intf_322(clock,reset);
    assign fifo_intf_322.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_14_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_14_U.if_empty_n;
    assign fifo_intf_322.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_14_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_14_U.if_full_n;
    assign fifo_intf_322.fifo_rd_block = 0;
    assign fifo_intf_322.fifo_wr_block = 0;
    assign fifo_intf_322.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_322;
    csv_file_dump cstatus_csv_dumper_322;
    df_fifo_monitor fifo_monitor_322;
    df_fifo_intf fifo_intf_323(clock,reset);
    assign fifo_intf_323.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_15_U.if_empty_n;
    assign fifo_intf_323.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_15_U.if_full_n;
    assign fifo_intf_323.fifo_rd_block = 0;
    assign fifo_intf_323.fifo_wr_block = 0;
    assign fifo_intf_323.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_323;
    csv_file_dump cstatus_csv_dumper_323;
    df_fifo_monitor fifo_monitor_323;
    df_fifo_intf fifo_intf_324(clock,reset);
    assign fifo_intf_324.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_15_U.if_empty_n;
    assign fifo_intf_324.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_15_U.if_full_n;
    assign fifo_intf_324.fifo_rd_block = 0;
    assign fifo_intf_324.fifo_wr_block = 0;
    assign fifo_intf_324.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_324;
    csv_file_dump cstatus_csv_dumper_324;
    df_fifo_monitor fifo_monitor_324;
    df_fifo_intf fifo_intf_325(clock,reset);
    assign fifo_intf_325.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_15_U.if_empty_n;
    assign fifo_intf_325.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_15_U.if_full_n;
    assign fifo_intf_325.fifo_rd_block = 0;
    assign fifo_intf_325.fifo_wr_block = 0;
    assign fifo_intf_325.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_325;
    csv_file_dump cstatus_csv_dumper_325;
    df_fifo_monitor fifo_monitor_325;
    df_fifo_intf fifo_intf_326(clock,reset);
    assign fifo_intf_326.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_15_U.if_empty_n;
    assign fifo_intf_326.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_15_U.if_full_n;
    assign fifo_intf_326.fifo_rd_block = 0;
    assign fifo_intf_326.fifo_wr_block = 0;
    assign fifo_intf_326.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_326;
    csv_file_dump cstatus_csv_dumper_326;
    df_fifo_monitor fifo_monitor_326;
    df_fifo_intf fifo_intf_327(clock,reset);
    assign fifo_intf_327.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_15_U.if_empty_n;
    assign fifo_intf_327.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_15_U.if_full_n;
    assign fifo_intf_327.fifo_rd_block = 0;
    assign fifo_intf_327.fifo_wr_block = 0;
    assign fifo_intf_327.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_327;
    csv_file_dump cstatus_csv_dumper_327;
    df_fifo_monitor fifo_monitor_327;
    df_fifo_intf fifo_intf_328(clock,reset);
    assign fifo_intf_328.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_15_U.if_empty_n;
    assign fifo_intf_328.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_15_U.if_full_n;
    assign fifo_intf_328.fifo_rd_block = 0;
    assign fifo_intf_328.fifo_wr_block = 0;
    assign fifo_intf_328.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_328;
    csv_file_dump cstatus_csv_dumper_328;
    df_fifo_monitor fifo_monitor_328;
    df_fifo_intf fifo_intf_329(clock,reset);
    assign fifo_intf_329.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_15_U.if_empty_n;
    assign fifo_intf_329.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_15_U.if_full_n;
    assign fifo_intf_329.fifo_rd_block = 0;
    assign fifo_intf_329.fifo_wr_block = 0;
    assign fifo_intf_329.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_329;
    csv_file_dump cstatus_csv_dumper_329;
    df_fifo_monitor fifo_monitor_329;
    df_fifo_intf fifo_intf_330(clock,reset);
    assign fifo_intf_330.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_15_U.if_empty_n;
    assign fifo_intf_330.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_15_U.if_full_n;
    assign fifo_intf_330.fifo_rd_block = 0;
    assign fifo_intf_330.fifo_wr_block = 0;
    assign fifo_intf_330.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_330;
    csv_file_dump cstatus_csv_dumper_330;
    df_fifo_monitor fifo_monitor_330;
    df_fifo_intf fifo_intf_331(clock,reset);
    assign fifo_intf_331.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_15_U.if_empty_n;
    assign fifo_intf_331.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_15_U.if_full_n;
    assign fifo_intf_331.fifo_rd_block = 0;
    assign fifo_intf_331.fifo_wr_block = 0;
    assign fifo_intf_331.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_331;
    csv_file_dump cstatus_csv_dumper_331;
    df_fifo_monitor fifo_monitor_331;
    df_fifo_intf fifo_intf_332(clock,reset);
    assign fifo_intf_332.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_15_U.if_empty_n;
    assign fifo_intf_332.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_15_U.if_full_n;
    assign fifo_intf_332.fifo_rd_block = 0;
    assign fifo_intf_332.fifo_wr_block = 0;
    assign fifo_intf_332.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_332;
    csv_file_dump cstatus_csv_dumper_332;
    df_fifo_monitor fifo_monitor_332;
    df_fifo_intf fifo_intf_333(clock,reset);
    assign fifo_intf_333.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_15_U.if_empty_n;
    assign fifo_intf_333.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_15_U.if_full_n;
    assign fifo_intf_333.fifo_rd_block = 0;
    assign fifo_intf_333.fifo_wr_block = 0;
    assign fifo_intf_333.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_333;
    csv_file_dump cstatus_csv_dumper_333;
    df_fifo_monitor fifo_monitor_333;
    df_fifo_intf fifo_intf_334(clock,reset);
    assign fifo_intf_334.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_15_U.if_empty_n;
    assign fifo_intf_334.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_15_U.if_full_n;
    assign fifo_intf_334.fifo_rd_block = 0;
    assign fifo_intf_334.fifo_wr_block = 0;
    assign fifo_intf_334.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_334;
    csv_file_dump cstatus_csv_dumper_334;
    df_fifo_monitor fifo_monitor_334;
    df_fifo_intf fifo_intf_335(clock,reset);
    assign fifo_intf_335.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_15_U.if_empty_n;
    assign fifo_intf_335.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_15_U.if_full_n;
    assign fifo_intf_335.fifo_rd_block = 0;
    assign fifo_intf_335.fifo_wr_block = 0;
    assign fifo_intf_335.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_335;
    csv_file_dump cstatus_csv_dumper_335;
    df_fifo_monitor fifo_monitor_335;
    df_fifo_intf fifo_intf_336(clock,reset);
    assign fifo_intf_336.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_15_U.if_empty_n;
    assign fifo_intf_336.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_15_U.if_full_n;
    assign fifo_intf_336.fifo_rd_block = 0;
    assign fifo_intf_336.fifo_wr_block = 0;
    assign fifo_intf_336.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_336;
    csv_file_dump cstatus_csv_dumper_336;
    df_fifo_monitor fifo_monitor_336;
    df_fifo_intf fifo_intf_337(clock,reset);
    assign fifo_intf_337.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_15_U.if_empty_n;
    assign fifo_intf_337.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_15_U.if_full_n;
    assign fifo_intf_337.fifo_rd_block = 0;
    assign fifo_intf_337.fifo_wr_block = 0;
    assign fifo_intf_337.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_337;
    csv_file_dump cstatus_csv_dumper_337;
    df_fifo_monitor fifo_monitor_337;
    df_fifo_intf fifo_intf_338(clock,reset);
    assign fifo_intf_338.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_15_U.if_empty_n;
    assign fifo_intf_338.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_15_U.if_full_n;
    assign fifo_intf_338.fifo_rd_block = 0;
    assign fifo_intf_338.fifo_wr_block = 0;
    assign fifo_intf_338.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_338;
    csv_file_dump cstatus_csv_dumper_338;
    df_fifo_monitor fifo_monitor_338;
    df_fifo_intf fifo_intf_339(clock,reset);
    assign fifo_intf_339.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_15_U.if_empty_n;
    assign fifo_intf_339.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_15_U.if_full_n;
    assign fifo_intf_339.fifo_rd_block = 0;
    assign fifo_intf_339.fifo_wr_block = 0;
    assign fifo_intf_339.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_339;
    csv_file_dump cstatus_csv_dumper_339;
    df_fifo_monitor fifo_monitor_339;
    df_fifo_intf fifo_intf_340(clock,reset);
    assign fifo_intf_340.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_15_U.if_empty_n;
    assign fifo_intf_340.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_15_U.if_full_n;
    assign fifo_intf_340.fifo_rd_block = 0;
    assign fifo_intf_340.fifo_wr_block = 0;
    assign fifo_intf_340.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_340;
    csv_file_dump cstatus_csv_dumper_340;
    df_fifo_monitor fifo_monitor_340;
    df_fifo_intf fifo_intf_341(clock,reset);
    assign fifo_intf_341.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_15_U.if_empty_n;
    assign fifo_intf_341.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_15_U.if_full_n;
    assign fifo_intf_341.fifo_rd_block = 0;
    assign fifo_intf_341.fifo_wr_block = 0;
    assign fifo_intf_341.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_341;
    csv_file_dump cstatus_csv_dumper_341;
    df_fifo_monitor fifo_monitor_341;
    df_fifo_intf fifo_intf_342(clock,reset);
    assign fifo_intf_342.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_15_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_15_U.if_empty_n;
    assign fifo_intf_342.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_15_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_15_U.if_full_n;
    assign fifo_intf_342.fifo_rd_block = 0;
    assign fifo_intf_342.fifo_wr_block = 0;
    assign fifo_intf_342.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_342;
    csv_file_dump cstatus_csv_dumper_342;
    df_fifo_monitor fifo_monitor_342;
    df_fifo_intf fifo_intf_343(clock,reset);
    assign fifo_intf_343.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_16_U.if_empty_n;
    assign fifo_intf_343.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_16_U.if_full_n;
    assign fifo_intf_343.fifo_rd_block = 0;
    assign fifo_intf_343.fifo_wr_block = 0;
    assign fifo_intf_343.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_343;
    csv_file_dump cstatus_csv_dumper_343;
    df_fifo_monitor fifo_monitor_343;
    df_fifo_intf fifo_intf_344(clock,reset);
    assign fifo_intf_344.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_16_U.if_empty_n;
    assign fifo_intf_344.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_16_U.if_full_n;
    assign fifo_intf_344.fifo_rd_block = 0;
    assign fifo_intf_344.fifo_wr_block = 0;
    assign fifo_intf_344.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_344;
    csv_file_dump cstatus_csv_dumper_344;
    df_fifo_monitor fifo_monitor_344;
    df_fifo_intf fifo_intf_345(clock,reset);
    assign fifo_intf_345.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_16_U.if_empty_n;
    assign fifo_intf_345.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_16_U.if_full_n;
    assign fifo_intf_345.fifo_rd_block = 0;
    assign fifo_intf_345.fifo_wr_block = 0;
    assign fifo_intf_345.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_345;
    csv_file_dump cstatus_csv_dumper_345;
    df_fifo_monitor fifo_monitor_345;
    df_fifo_intf fifo_intf_346(clock,reset);
    assign fifo_intf_346.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_16_U.if_empty_n;
    assign fifo_intf_346.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_16_U.if_full_n;
    assign fifo_intf_346.fifo_rd_block = 0;
    assign fifo_intf_346.fifo_wr_block = 0;
    assign fifo_intf_346.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_346;
    csv_file_dump cstatus_csv_dumper_346;
    df_fifo_monitor fifo_monitor_346;
    df_fifo_intf fifo_intf_347(clock,reset);
    assign fifo_intf_347.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_16_U.if_empty_n;
    assign fifo_intf_347.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_16_U.if_full_n;
    assign fifo_intf_347.fifo_rd_block = 0;
    assign fifo_intf_347.fifo_wr_block = 0;
    assign fifo_intf_347.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_347;
    csv_file_dump cstatus_csv_dumper_347;
    df_fifo_monitor fifo_monitor_347;
    df_fifo_intf fifo_intf_348(clock,reset);
    assign fifo_intf_348.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_16_U.if_empty_n;
    assign fifo_intf_348.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_16_U.if_full_n;
    assign fifo_intf_348.fifo_rd_block = 0;
    assign fifo_intf_348.fifo_wr_block = 0;
    assign fifo_intf_348.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_348;
    csv_file_dump cstatus_csv_dumper_348;
    df_fifo_monitor fifo_monitor_348;
    df_fifo_intf fifo_intf_349(clock,reset);
    assign fifo_intf_349.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_16_U.if_empty_n;
    assign fifo_intf_349.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_16_U.if_full_n;
    assign fifo_intf_349.fifo_rd_block = 0;
    assign fifo_intf_349.fifo_wr_block = 0;
    assign fifo_intf_349.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_349;
    csv_file_dump cstatus_csv_dumper_349;
    df_fifo_monitor fifo_monitor_349;
    df_fifo_intf fifo_intf_350(clock,reset);
    assign fifo_intf_350.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_16_U.if_empty_n;
    assign fifo_intf_350.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_16_U.if_full_n;
    assign fifo_intf_350.fifo_rd_block = 0;
    assign fifo_intf_350.fifo_wr_block = 0;
    assign fifo_intf_350.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_350;
    csv_file_dump cstatus_csv_dumper_350;
    df_fifo_monitor fifo_monitor_350;
    df_fifo_intf fifo_intf_351(clock,reset);
    assign fifo_intf_351.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_16_U.if_empty_n;
    assign fifo_intf_351.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_16_U.if_full_n;
    assign fifo_intf_351.fifo_rd_block = 0;
    assign fifo_intf_351.fifo_wr_block = 0;
    assign fifo_intf_351.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_351;
    csv_file_dump cstatus_csv_dumper_351;
    df_fifo_monitor fifo_monitor_351;
    df_fifo_intf fifo_intf_352(clock,reset);
    assign fifo_intf_352.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_16_U.if_empty_n;
    assign fifo_intf_352.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_16_U.if_full_n;
    assign fifo_intf_352.fifo_rd_block = 0;
    assign fifo_intf_352.fifo_wr_block = 0;
    assign fifo_intf_352.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_352;
    csv_file_dump cstatus_csv_dumper_352;
    df_fifo_monitor fifo_monitor_352;
    df_fifo_intf fifo_intf_353(clock,reset);
    assign fifo_intf_353.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_16_U.if_empty_n;
    assign fifo_intf_353.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_16_U.if_full_n;
    assign fifo_intf_353.fifo_rd_block = 0;
    assign fifo_intf_353.fifo_wr_block = 0;
    assign fifo_intf_353.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_353;
    csv_file_dump cstatus_csv_dumper_353;
    df_fifo_monitor fifo_monitor_353;
    df_fifo_intf fifo_intf_354(clock,reset);
    assign fifo_intf_354.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_16_U.if_empty_n;
    assign fifo_intf_354.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_16_U.if_full_n;
    assign fifo_intf_354.fifo_rd_block = 0;
    assign fifo_intf_354.fifo_wr_block = 0;
    assign fifo_intf_354.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_354;
    csv_file_dump cstatus_csv_dumper_354;
    df_fifo_monitor fifo_monitor_354;
    df_fifo_intf fifo_intf_355(clock,reset);
    assign fifo_intf_355.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_16_U.if_empty_n;
    assign fifo_intf_355.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_16_U.if_full_n;
    assign fifo_intf_355.fifo_rd_block = 0;
    assign fifo_intf_355.fifo_wr_block = 0;
    assign fifo_intf_355.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_355;
    csv_file_dump cstatus_csv_dumper_355;
    df_fifo_monitor fifo_monitor_355;
    df_fifo_intf fifo_intf_356(clock,reset);
    assign fifo_intf_356.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_16_U.if_empty_n;
    assign fifo_intf_356.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_16_U.if_full_n;
    assign fifo_intf_356.fifo_rd_block = 0;
    assign fifo_intf_356.fifo_wr_block = 0;
    assign fifo_intf_356.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_356;
    csv_file_dump cstatus_csv_dumper_356;
    df_fifo_monitor fifo_monitor_356;
    df_fifo_intf fifo_intf_357(clock,reset);
    assign fifo_intf_357.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_16_U.if_empty_n;
    assign fifo_intf_357.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_16_U.if_full_n;
    assign fifo_intf_357.fifo_rd_block = 0;
    assign fifo_intf_357.fifo_wr_block = 0;
    assign fifo_intf_357.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_357;
    csv_file_dump cstatus_csv_dumper_357;
    df_fifo_monitor fifo_monitor_357;
    df_fifo_intf fifo_intf_358(clock,reset);
    assign fifo_intf_358.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_16_U.if_empty_n;
    assign fifo_intf_358.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_16_U.if_full_n;
    assign fifo_intf_358.fifo_rd_block = 0;
    assign fifo_intf_358.fifo_wr_block = 0;
    assign fifo_intf_358.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_358;
    csv_file_dump cstatus_csv_dumper_358;
    df_fifo_monitor fifo_monitor_358;
    df_fifo_intf fifo_intf_359(clock,reset);
    assign fifo_intf_359.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_16_U.if_empty_n;
    assign fifo_intf_359.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_16_U.if_full_n;
    assign fifo_intf_359.fifo_rd_block = 0;
    assign fifo_intf_359.fifo_wr_block = 0;
    assign fifo_intf_359.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_359;
    csv_file_dump cstatus_csv_dumper_359;
    df_fifo_monitor fifo_monitor_359;
    df_fifo_intf fifo_intf_360(clock,reset);
    assign fifo_intf_360.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_16_U.if_empty_n;
    assign fifo_intf_360.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_16_U.if_full_n;
    assign fifo_intf_360.fifo_rd_block = 0;
    assign fifo_intf_360.fifo_wr_block = 0;
    assign fifo_intf_360.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_360;
    csv_file_dump cstatus_csv_dumper_360;
    df_fifo_monitor fifo_monitor_360;
    df_fifo_intf fifo_intf_361(clock,reset);
    assign fifo_intf_361.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_16_U.if_empty_n;
    assign fifo_intf_361.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_16_U.if_full_n;
    assign fifo_intf_361.fifo_rd_block = 0;
    assign fifo_intf_361.fifo_wr_block = 0;
    assign fifo_intf_361.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_361;
    csv_file_dump cstatus_csv_dumper_361;
    df_fifo_monitor fifo_monitor_361;
    df_fifo_intf fifo_intf_362(clock,reset);
    assign fifo_intf_362.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_16_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_16_U.if_empty_n;
    assign fifo_intf_362.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_16_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_16_U.if_full_n;
    assign fifo_intf_362.fifo_rd_block = 0;
    assign fifo_intf_362.fifo_wr_block = 0;
    assign fifo_intf_362.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_362;
    csv_file_dump cstatus_csv_dumper_362;
    df_fifo_monitor fifo_monitor_362;
    df_fifo_intf fifo_intf_363(clock,reset);
    assign fifo_intf_363.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_17_U.if_empty_n;
    assign fifo_intf_363.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_17_U.if_full_n;
    assign fifo_intf_363.fifo_rd_block = 0;
    assign fifo_intf_363.fifo_wr_block = 0;
    assign fifo_intf_363.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_363;
    csv_file_dump cstatus_csv_dumper_363;
    df_fifo_monitor fifo_monitor_363;
    df_fifo_intf fifo_intf_364(clock,reset);
    assign fifo_intf_364.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_17_U.if_empty_n;
    assign fifo_intf_364.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_17_U.if_full_n;
    assign fifo_intf_364.fifo_rd_block = 0;
    assign fifo_intf_364.fifo_wr_block = 0;
    assign fifo_intf_364.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_364;
    csv_file_dump cstatus_csv_dumper_364;
    df_fifo_monitor fifo_monitor_364;
    df_fifo_intf fifo_intf_365(clock,reset);
    assign fifo_intf_365.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_17_U.if_empty_n;
    assign fifo_intf_365.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_17_U.if_full_n;
    assign fifo_intf_365.fifo_rd_block = 0;
    assign fifo_intf_365.fifo_wr_block = 0;
    assign fifo_intf_365.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_365;
    csv_file_dump cstatus_csv_dumper_365;
    df_fifo_monitor fifo_monitor_365;
    df_fifo_intf fifo_intf_366(clock,reset);
    assign fifo_intf_366.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_17_U.if_empty_n;
    assign fifo_intf_366.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_17_U.if_full_n;
    assign fifo_intf_366.fifo_rd_block = 0;
    assign fifo_intf_366.fifo_wr_block = 0;
    assign fifo_intf_366.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_366;
    csv_file_dump cstatus_csv_dumper_366;
    df_fifo_monitor fifo_monitor_366;
    df_fifo_intf fifo_intf_367(clock,reset);
    assign fifo_intf_367.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_17_U.if_empty_n;
    assign fifo_intf_367.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_17_U.if_full_n;
    assign fifo_intf_367.fifo_rd_block = 0;
    assign fifo_intf_367.fifo_wr_block = 0;
    assign fifo_intf_367.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_367;
    csv_file_dump cstatus_csv_dumper_367;
    df_fifo_monitor fifo_monitor_367;
    df_fifo_intf fifo_intf_368(clock,reset);
    assign fifo_intf_368.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_17_U.if_empty_n;
    assign fifo_intf_368.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_17_U.if_full_n;
    assign fifo_intf_368.fifo_rd_block = 0;
    assign fifo_intf_368.fifo_wr_block = 0;
    assign fifo_intf_368.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_368;
    csv_file_dump cstatus_csv_dumper_368;
    df_fifo_monitor fifo_monitor_368;
    df_fifo_intf fifo_intf_369(clock,reset);
    assign fifo_intf_369.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_17_U.if_empty_n;
    assign fifo_intf_369.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_17_U.if_full_n;
    assign fifo_intf_369.fifo_rd_block = 0;
    assign fifo_intf_369.fifo_wr_block = 0;
    assign fifo_intf_369.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_369;
    csv_file_dump cstatus_csv_dumper_369;
    df_fifo_monitor fifo_monitor_369;
    df_fifo_intf fifo_intf_370(clock,reset);
    assign fifo_intf_370.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_17_U.if_empty_n;
    assign fifo_intf_370.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_17_U.if_full_n;
    assign fifo_intf_370.fifo_rd_block = 0;
    assign fifo_intf_370.fifo_wr_block = 0;
    assign fifo_intf_370.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_370;
    csv_file_dump cstatus_csv_dumper_370;
    df_fifo_monitor fifo_monitor_370;
    df_fifo_intf fifo_intf_371(clock,reset);
    assign fifo_intf_371.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_17_U.if_empty_n;
    assign fifo_intf_371.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_17_U.if_full_n;
    assign fifo_intf_371.fifo_rd_block = 0;
    assign fifo_intf_371.fifo_wr_block = 0;
    assign fifo_intf_371.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_371;
    csv_file_dump cstatus_csv_dumper_371;
    df_fifo_monitor fifo_monitor_371;
    df_fifo_intf fifo_intf_372(clock,reset);
    assign fifo_intf_372.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_17_U.if_empty_n;
    assign fifo_intf_372.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_17_U.if_full_n;
    assign fifo_intf_372.fifo_rd_block = 0;
    assign fifo_intf_372.fifo_wr_block = 0;
    assign fifo_intf_372.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_372;
    csv_file_dump cstatus_csv_dumper_372;
    df_fifo_monitor fifo_monitor_372;
    df_fifo_intf fifo_intf_373(clock,reset);
    assign fifo_intf_373.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_17_U.if_empty_n;
    assign fifo_intf_373.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_17_U.if_full_n;
    assign fifo_intf_373.fifo_rd_block = 0;
    assign fifo_intf_373.fifo_wr_block = 0;
    assign fifo_intf_373.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_373;
    csv_file_dump cstatus_csv_dumper_373;
    df_fifo_monitor fifo_monitor_373;
    df_fifo_intf fifo_intf_374(clock,reset);
    assign fifo_intf_374.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_17_U.if_empty_n;
    assign fifo_intf_374.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_17_U.if_full_n;
    assign fifo_intf_374.fifo_rd_block = 0;
    assign fifo_intf_374.fifo_wr_block = 0;
    assign fifo_intf_374.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_374;
    csv_file_dump cstatus_csv_dumper_374;
    df_fifo_monitor fifo_monitor_374;
    df_fifo_intf fifo_intf_375(clock,reset);
    assign fifo_intf_375.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_17_U.if_empty_n;
    assign fifo_intf_375.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_17_U.if_full_n;
    assign fifo_intf_375.fifo_rd_block = 0;
    assign fifo_intf_375.fifo_wr_block = 0;
    assign fifo_intf_375.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_375;
    csv_file_dump cstatus_csv_dumper_375;
    df_fifo_monitor fifo_monitor_375;
    df_fifo_intf fifo_intf_376(clock,reset);
    assign fifo_intf_376.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_17_U.if_empty_n;
    assign fifo_intf_376.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_17_U.if_full_n;
    assign fifo_intf_376.fifo_rd_block = 0;
    assign fifo_intf_376.fifo_wr_block = 0;
    assign fifo_intf_376.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_376;
    csv_file_dump cstatus_csv_dumper_376;
    df_fifo_monitor fifo_monitor_376;
    df_fifo_intf fifo_intf_377(clock,reset);
    assign fifo_intf_377.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_17_U.if_empty_n;
    assign fifo_intf_377.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_17_U.if_full_n;
    assign fifo_intf_377.fifo_rd_block = 0;
    assign fifo_intf_377.fifo_wr_block = 0;
    assign fifo_intf_377.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_377;
    csv_file_dump cstatus_csv_dumper_377;
    df_fifo_monitor fifo_monitor_377;
    df_fifo_intf fifo_intf_378(clock,reset);
    assign fifo_intf_378.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_17_U.if_empty_n;
    assign fifo_intf_378.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_17_U.if_full_n;
    assign fifo_intf_378.fifo_rd_block = 0;
    assign fifo_intf_378.fifo_wr_block = 0;
    assign fifo_intf_378.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_378;
    csv_file_dump cstatus_csv_dumper_378;
    df_fifo_monitor fifo_monitor_378;
    df_fifo_intf fifo_intf_379(clock,reset);
    assign fifo_intf_379.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_17_U.if_empty_n;
    assign fifo_intf_379.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_17_U.if_full_n;
    assign fifo_intf_379.fifo_rd_block = 0;
    assign fifo_intf_379.fifo_wr_block = 0;
    assign fifo_intf_379.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_379;
    csv_file_dump cstatus_csv_dumper_379;
    df_fifo_monitor fifo_monitor_379;
    df_fifo_intf fifo_intf_380(clock,reset);
    assign fifo_intf_380.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_17_U.if_empty_n;
    assign fifo_intf_380.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_17_U.if_full_n;
    assign fifo_intf_380.fifo_rd_block = 0;
    assign fifo_intf_380.fifo_wr_block = 0;
    assign fifo_intf_380.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_380;
    csv_file_dump cstatus_csv_dumper_380;
    df_fifo_monitor fifo_monitor_380;
    df_fifo_intf fifo_intf_381(clock,reset);
    assign fifo_intf_381.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_17_U.if_empty_n;
    assign fifo_intf_381.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_17_U.if_full_n;
    assign fifo_intf_381.fifo_rd_block = 0;
    assign fifo_intf_381.fifo_wr_block = 0;
    assign fifo_intf_381.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_381;
    csv_file_dump cstatus_csv_dumper_381;
    df_fifo_monitor fifo_monitor_381;
    df_fifo_intf fifo_intf_382(clock,reset);
    assign fifo_intf_382.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_17_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_17_U.if_empty_n;
    assign fifo_intf_382.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_17_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_17_U.if_full_n;
    assign fifo_intf_382.fifo_rd_block = 0;
    assign fifo_intf_382.fifo_wr_block = 0;
    assign fifo_intf_382.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_382;
    csv_file_dump cstatus_csv_dumper_382;
    df_fifo_monitor fifo_monitor_382;
    df_fifo_intf fifo_intf_383(clock,reset);
    assign fifo_intf_383.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_18_U.if_empty_n;
    assign fifo_intf_383.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_18_U.if_full_n;
    assign fifo_intf_383.fifo_rd_block = 0;
    assign fifo_intf_383.fifo_wr_block = 0;
    assign fifo_intf_383.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_383;
    csv_file_dump cstatus_csv_dumper_383;
    df_fifo_monitor fifo_monitor_383;
    df_fifo_intf fifo_intf_384(clock,reset);
    assign fifo_intf_384.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_18_U.if_empty_n;
    assign fifo_intf_384.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_18_U.if_full_n;
    assign fifo_intf_384.fifo_rd_block = 0;
    assign fifo_intf_384.fifo_wr_block = 0;
    assign fifo_intf_384.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_384;
    csv_file_dump cstatus_csv_dumper_384;
    df_fifo_monitor fifo_monitor_384;
    df_fifo_intf fifo_intf_385(clock,reset);
    assign fifo_intf_385.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_18_U.if_empty_n;
    assign fifo_intf_385.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_18_U.if_full_n;
    assign fifo_intf_385.fifo_rd_block = 0;
    assign fifo_intf_385.fifo_wr_block = 0;
    assign fifo_intf_385.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_385;
    csv_file_dump cstatus_csv_dumper_385;
    df_fifo_monitor fifo_monitor_385;
    df_fifo_intf fifo_intf_386(clock,reset);
    assign fifo_intf_386.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_18_U.if_empty_n;
    assign fifo_intf_386.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_18_U.if_full_n;
    assign fifo_intf_386.fifo_rd_block = 0;
    assign fifo_intf_386.fifo_wr_block = 0;
    assign fifo_intf_386.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_386;
    csv_file_dump cstatus_csv_dumper_386;
    df_fifo_monitor fifo_monitor_386;
    df_fifo_intf fifo_intf_387(clock,reset);
    assign fifo_intf_387.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_18_U.if_empty_n;
    assign fifo_intf_387.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_18_U.if_full_n;
    assign fifo_intf_387.fifo_rd_block = 0;
    assign fifo_intf_387.fifo_wr_block = 0;
    assign fifo_intf_387.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_387;
    csv_file_dump cstatus_csv_dumper_387;
    df_fifo_monitor fifo_monitor_387;
    df_fifo_intf fifo_intf_388(clock,reset);
    assign fifo_intf_388.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_18_U.if_empty_n;
    assign fifo_intf_388.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_18_U.if_full_n;
    assign fifo_intf_388.fifo_rd_block = 0;
    assign fifo_intf_388.fifo_wr_block = 0;
    assign fifo_intf_388.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_388;
    csv_file_dump cstatus_csv_dumper_388;
    df_fifo_monitor fifo_monitor_388;
    df_fifo_intf fifo_intf_389(clock,reset);
    assign fifo_intf_389.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_18_U.if_empty_n;
    assign fifo_intf_389.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_18_U.if_full_n;
    assign fifo_intf_389.fifo_rd_block = 0;
    assign fifo_intf_389.fifo_wr_block = 0;
    assign fifo_intf_389.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_389;
    csv_file_dump cstatus_csv_dumper_389;
    df_fifo_monitor fifo_monitor_389;
    df_fifo_intf fifo_intf_390(clock,reset);
    assign fifo_intf_390.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_18_U.if_empty_n;
    assign fifo_intf_390.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_18_U.if_full_n;
    assign fifo_intf_390.fifo_rd_block = 0;
    assign fifo_intf_390.fifo_wr_block = 0;
    assign fifo_intf_390.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_390;
    csv_file_dump cstatus_csv_dumper_390;
    df_fifo_monitor fifo_monitor_390;
    df_fifo_intf fifo_intf_391(clock,reset);
    assign fifo_intf_391.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_18_U.if_empty_n;
    assign fifo_intf_391.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_18_U.if_full_n;
    assign fifo_intf_391.fifo_rd_block = 0;
    assign fifo_intf_391.fifo_wr_block = 0;
    assign fifo_intf_391.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_391;
    csv_file_dump cstatus_csv_dumper_391;
    df_fifo_monitor fifo_monitor_391;
    df_fifo_intf fifo_intf_392(clock,reset);
    assign fifo_intf_392.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_18_U.if_empty_n;
    assign fifo_intf_392.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_18_U.if_full_n;
    assign fifo_intf_392.fifo_rd_block = 0;
    assign fifo_intf_392.fifo_wr_block = 0;
    assign fifo_intf_392.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_392;
    csv_file_dump cstatus_csv_dumper_392;
    df_fifo_monitor fifo_monitor_392;
    df_fifo_intf fifo_intf_393(clock,reset);
    assign fifo_intf_393.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_18_U.if_empty_n;
    assign fifo_intf_393.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_18_U.if_full_n;
    assign fifo_intf_393.fifo_rd_block = 0;
    assign fifo_intf_393.fifo_wr_block = 0;
    assign fifo_intf_393.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_393;
    csv_file_dump cstatus_csv_dumper_393;
    df_fifo_monitor fifo_monitor_393;
    df_fifo_intf fifo_intf_394(clock,reset);
    assign fifo_intf_394.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_18_U.if_empty_n;
    assign fifo_intf_394.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_18_U.if_full_n;
    assign fifo_intf_394.fifo_rd_block = 0;
    assign fifo_intf_394.fifo_wr_block = 0;
    assign fifo_intf_394.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_394;
    csv_file_dump cstatus_csv_dumper_394;
    df_fifo_monitor fifo_monitor_394;
    df_fifo_intf fifo_intf_395(clock,reset);
    assign fifo_intf_395.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_18_U.if_empty_n;
    assign fifo_intf_395.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_18_U.if_full_n;
    assign fifo_intf_395.fifo_rd_block = 0;
    assign fifo_intf_395.fifo_wr_block = 0;
    assign fifo_intf_395.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_395;
    csv_file_dump cstatus_csv_dumper_395;
    df_fifo_monitor fifo_monitor_395;
    df_fifo_intf fifo_intf_396(clock,reset);
    assign fifo_intf_396.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_18_U.if_empty_n;
    assign fifo_intf_396.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_18_U.if_full_n;
    assign fifo_intf_396.fifo_rd_block = 0;
    assign fifo_intf_396.fifo_wr_block = 0;
    assign fifo_intf_396.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_396;
    csv_file_dump cstatus_csv_dumper_396;
    df_fifo_monitor fifo_monitor_396;
    df_fifo_intf fifo_intf_397(clock,reset);
    assign fifo_intf_397.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_18_U.if_empty_n;
    assign fifo_intf_397.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_18_U.if_full_n;
    assign fifo_intf_397.fifo_rd_block = 0;
    assign fifo_intf_397.fifo_wr_block = 0;
    assign fifo_intf_397.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_397;
    csv_file_dump cstatus_csv_dumper_397;
    df_fifo_monitor fifo_monitor_397;
    df_fifo_intf fifo_intf_398(clock,reset);
    assign fifo_intf_398.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_18_U.if_empty_n;
    assign fifo_intf_398.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_18_U.if_full_n;
    assign fifo_intf_398.fifo_rd_block = 0;
    assign fifo_intf_398.fifo_wr_block = 0;
    assign fifo_intf_398.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_398;
    csv_file_dump cstatus_csv_dumper_398;
    df_fifo_monitor fifo_monitor_398;
    df_fifo_intf fifo_intf_399(clock,reset);
    assign fifo_intf_399.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_18_U.if_empty_n;
    assign fifo_intf_399.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_18_U.if_full_n;
    assign fifo_intf_399.fifo_rd_block = 0;
    assign fifo_intf_399.fifo_wr_block = 0;
    assign fifo_intf_399.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_399;
    csv_file_dump cstatus_csv_dumper_399;
    df_fifo_monitor fifo_monitor_399;
    df_fifo_intf fifo_intf_400(clock,reset);
    assign fifo_intf_400.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_18_U.if_empty_n;
    assign fifo_intf_400.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_18_U.if_full_n;
    assign fifo_intf_400.fifo_rd_block = 0;
    assign fifo_intf_400.fifo_wr_block = 0;
    assign fifo_intf_400.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_400;
    csv_file_dump cstatus_csv_dumper_400;
    df_fifo_monitor fifo_monitor_400;
    df_fifo_intf fifo_intf_401(clock,reset);
    assign fifo_intf_401.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_18_U.if_empty_n;
    assign fifo_intf_401.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_18_U.if_full_n;
    assign fifo_intf_401.fifo_rd_block = 0;
    assign fifo_intf_401.fifo_wr_block = 0;
    assign fifo_intf_401.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_401;
    csv_file_dump cstatus_csv_dumper_401;
    df_fifo_monitor fifo_monitor_401;
    df_fifo_intf fifo_intf_402(clock,reset);
    assign fifo_intf_402.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_18_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_18_U.if_empty_n;
    assign fifo_intf_402.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_18_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_18_U.if_full_n;
    assign fifo_intf_402.fifo_rd_block = 0;
    assign fifo_intf_402.fifo_wr_block = 0;
    assign fifo_intf_402.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_402;
    csv_file_dump cstatus_csv_dumper_402;
    df_fifo_monitor fifo_monitor_402;
    df_fifo_intf fifo_intf_403(clock,reset);
    assign fifo_intf_403.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_19_U.if_empty_n;
    assign fifo_intf_403.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_19_U.if_full_n;
    assign fifo_intf_403.fifo_rd_block = 0;
    assign fifo_intf_403.fifo_wr_block = 0;
    assign fifo_intf_403.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_403;
    csv_file_dump cstatus_csv_dumper_403;
    df_fifo_monitor fifo_monitor_403;
    df_fifo_intf fifo_intf_404(clock,reset);
    assign fifo_intf_404.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_19_U.if_empty_n;
    assign fifo_intf_404.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_19_U.if_full_n;
    assign fifo_intf_404.fifo_rd_block = 0;
    assign fifo_intf_404.fifo_wr_block = 0;
    assign fifo_intf_404.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_404;
    csv_file_dump cstatus_csv_dumper_404;
    df_fifo_monitor fifo_monitor_404;
    df_fifo_intf fifo_intf_405(clock,reset);
    assign fifo_intf_405.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_19_U.if_empty_n;
    assign fifo_intf_405.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_19_U.if_full_n;
    assign fifo_intf_405.fifo_rd_block = 0;
    assign fifo_intf_405.fifo_wr_block = 0;
    assign fifo_intf_405.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_405;
    csv_file_dump cstatus_csv_dumper_405;
    df_fifo_monitor fifo_monitor_405;
    df_fifo_intf fifo_intf_406(clock,reset);
    assign fifo_intf_406.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_19_U.if_empty_n;
    assign fifo_intf_406.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_19_U.if_full_n;
    assign fifo_intf_406.fifo_rd_block = 0;
    assign fifo_intf_406.fifo_wr_block = 0;
    assign fifo_intf_406.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_406;
    csv_file_dump cstatus_csv_dumper_406;
    df_fifo_monitor fifo_monitor_406;
    df_fifo_intf fifo_intf_407(clock,reset);
    assign fifo_intf_407.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_19_U.if_empty_n;
    assign fifo_intf_407.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_19_U.if_full_n;
    assign fifo_intf_407.fifo_rd_block = 0;
    assign fifo_intf_407.fifo_wr_block = 0;
    assign fifo_intf_407.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_407;
    csv_file_dump cstatus_csv_dumper_407;
    df_fifo_monitor fifo_monitor_407;
    df_fifo_intf fifo_intf_408(clock,reset);
    assign fifo_intf_408.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_19_U.if_empty_n;
    assign fifo_intf_408.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_19_U.if_full_n;
    assign fifo_intf_408.fifo_rd_block = 0;
    assign fifo_intf_408.fifo_wr_block = 0;
    assign fifo_intf_408.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_408;
    csv_file_dump cstatus_csv_dumper_408;
    df_fifo_monitor fifo_monitor_408;
    df_fifo_intf fifo_intf_409(clock,reset);
    assign fifo_intf_409.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_19_U.if_empty_n;
    assign fifo_intf_409.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_19_U.if_full_n;
    assign fifo_intf_409.fifo_rd_block = 0;
    assign fifo_intf_409.fifo_wr_block = 0;
    assign fifo_intf_409.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_409;
    csv_file_dump cstatus_csv_dumper_409;
    df_fifo_monitor fifo_monitor_409;
    df_fifo_intf fifo_intf_410(clock,reset);
    assign fifo_intf_410.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_19_U.if_empty_n;
    assign fifo_intf_410.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_19_U.if_full_n;
    assign fifo_intf_410.fifo_rd_block = 0;
    assign fifo_intf_410.fifo_wr_block = 0;
    assign fifo_intf_410.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_410;
    csv_file_dump cstatus_csv_dumper_410;
    df_fifo_monitor fifo_monitor_410;
    df_fifo_intf fifo_intf_411(clock,reset);
    assign fifo_intf_411.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_19_U.if_empty_n;
    assign fifo_intf_411.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_19_U.if_full_n;
    assign fifo_intf_411.fifo_rd_block = 0;
    assign fifo_intf_411.fifo_wr_block = 0;
    assign fifo_intf_411.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_411;
    csv_file_dump cstatus_csv_dumper_411;
    df_fifo_monitor fifo_monitor_411;
    df_fifo_intf fifo_intf_412(clock,reset);
    assign fifo_intf_412.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_19_U.if_empty_n;
    assign fifo_intf_412.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_19_U.if_full_n;
    assign fifo_intf_412.fifo_rd_block = 0;
    assign fifo_intf_412.fifo_wr_block = 0;
    assign fifo_intf_412.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_412;
    csv_file_dump cstatus_csv_dumper_412;
    df_fifo_monitor fifo_monitor_412;
    df_fifo_intf fifo_intf_413(clock,reset);
    assign fifo_intf_413.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_19_U.if_empty_n;
    assign fifo_intf_413.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_19_U.if_full_n;
    assign fifo_intf_413.fifo_rd_block = 0;
    assign fifo_intf_413.fifo_wr_block = 0;
    assign fifo_intf_413.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_413;
    csv_file_dump cstatus_csv_dumper_413;
    df_fifo_monitor fifo_monitor_413;
    df_fifo_intf fifo_intf_414(clock,reset);
    assign fifo_intf_414.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_19_U.if_empty_n;
    assign fifo_intf_414.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_19_U.if_full_n;
    assign fifo_intf_414.fifo_rd_block = 0;
    assign fifo_intf_414.fifo_wr_block = 0;
    assign fifo_intf_414.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_414;
    csv_file_dump cstatus_csv_dumper_414;
    df_fifo_monitor fifo_monitor_414;
    df_fifo_intf fifo_intf_415(clock,reset);
    assign fifo_intf_415.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_19_U.if_empty_n;
    assign fifo_intf_415.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_19_U.if_full_n;
    assign fifo_intf_415.fifo_rd_block = 0;
    assign fifo_intf_415.fifo_wr_block = 0;
    assign fifo_intf_415.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_415;
    csv_file_dump cstatus_csv_dumper_415;
    df_fifo_monitor fifo_monitor_415;
    df_fifo_intf fifo_intf_416(clock,reset);
    assign fifo_intf_416.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_19_U.if_empty_n;
    assign fifo_intf_416.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_19_U.if_full_n;
    assign fifo_intf_416.fifo_rd_block = 0;
    assign fifo_intf_416.fifo_wr_block = 0;
    assign fifo_intf_416.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_416;
    csv_file_dump cstatus_csv_dumper_416;
    df_fifo_monitor fifo_monitor_416;
    df_fifo_intf fifo_intf_417(clock,reset);
    assign fifo_intf_417.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_19_U.if_empty_n;
    assign fifo_intf_417.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_19_U.if_full_n;
    assign fifo_intf_417.fifo_rd_block = 0;
    assign fifo_intf_417.fifo_wr_block = 0;
    assign fifo_intf_417.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_417;
    csv_file_dump cstatus_csv_dumper_417;
    df_fifo_monitor fifo_monitor_417;
    df_fifo_intf fifo_intf_418(clock,reset);
    assign fifo_intf_418.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_19_U.if_empty_n;
    assign fifo_intf_418.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_19_U.if_full_n;
    assign fifo_intf_418.fifo_rd_block = 0;
    assign fifo_intf_418.fifo_wr_block = 0;
    assign fifo_intf_418.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_418;
    csv_file_dump cstatus_csv_dumper_418;
    df_fifo_monitor fifo_monitor_418;
    df_fifo_intf fifo_intf_419(clock,reset);
    assign fifo_intf_419.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_19_U.if_empty_n;
    assign fifo_intf_419.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_19_U.if_full_n;
    assign fifo_intf_419.fifo_rd_block = 0;
    assign fifo_intf_419.fifo_wr_block = 0;
    assign fifo_intf_419.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_419;
    csv_file_dump cstatus_csv_dumper_419;
    df_fifo_monitor fifo_monitor_419;
    df_fifo_intf fifo_intf_420(clock,reset);
    assign fifo_intf_420.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_19_U.if_empty_n;
    assign fifo_intf_420.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_19_U.if_full_n;
    assign fifo_intf_420.fifo_rd_block = 0;
    assign fifo_intf_420.fifo_wr_block = 0;
    assign fifo_intf_420.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_420;
    csv_file_dump cstatus_csv_dumper_420;
    df_fifo_monitor fifo_monitor_420;
    df_fifo_intf fifo_intf_421(clock,reset);
    assign fifo_intf_421.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_19_U.if_empty_n;
    assign fifo_intf_421.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_19_U.if_full_n;
    assign fifo_intf_421.fifo_rd_block = 0;
    assign fifo_intf_421.fifo_wr_block = 0;
    assign fifo_intf_421.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_421;
    csv_file_dump cstatus_csv_dumper_421;
    df_fifo_monitor fifo_monitor_421;
    df_fifo_intf fifo_intf_422(clock,reset);
    assign fifo_intf_422.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_19_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_19_U.if_empty_n;
    assign fifo_intf_422.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_19_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_19_U.if_full_n;
    assign fifo_intf_422.fifo_rd_block = 0;
    assign fifo_intf_422.fifo_wr_block = 0;
    assign fifo_intf_422.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_422;
    csv_file_dump cstatus_csv_dumper_422;
    df_fifo_monitor fifo_monitor_422;
    df_fifo_intf fifo_intf_423(clock,reset);
    assign fifo_intf_423.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_U.if_empty_n;
    assign fifo_intf_423.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_U.if_full_n;
    assign fifo_intf_423.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_0_0_blk_n);
    assign fifo_intf_423.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.matr_out_0_0_blk_n);
    assign fifo_intf_423.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_423;
    csv_file_dump cstatus_csv_dumper_423;
    df_fifo_monitor fifo_monitor_423;
    df_fifo_intf fifo_intf_424(clock,reset);
    assign fifo_intf_424.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_1_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_1_U.if_empty_n;
    assign fifo_intf_424.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_1_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_1_U.if_full_n;
    assign fifo_intf_424.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_0_1_blk_n);
    assign fifo_intf_424.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.matr_out_0_1_blk_n);
    assign fifo_intf_424.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_424;
    csv_file_dump cstatus_csv_dumper_424;
    df_fifo_monitor fifo_monitor_424;
    df_fifo_intf fifo_intf_425(clock,reset);
    assign fifo_intf_425.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_20_U.if_empty_n;
    assign fifo_intf_425.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_20_U.if_full_n;
    assign fifo_intf_425.fifo_rd_block = 0;
    assign fifo_intf_425.fifo_wr_block = 0;
    assign fifo_intf_425.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_425;
    csv_file_dump cstatus_csv_dumper_425;
    df_fifo_monitor fifo_monitor_425;
    df_fifo_intf fifo_intf_426(clock,reset);
    assign fifo_intf_426.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_20_U.if_empty_n;
    assign fifo_intf_426.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_20_U.if_full_n;
    assign fifo_intf_426.fifo_rd_block = 0;
    assign fifo_intf_426.fifo_wr_block = 0;
    assign fifo_intf_426.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_426;
    csv_file_dump cstatus_csv_dumper_426;
    df_fifo_monitor fifo_monitor_426;
    df_fifo_intf fifo_intf_427(clock,reset);
    assign fifo_intf_427.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_20_U.if_empty_n;
    assign fifo_intf_427.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_20_U.if_full_n;
    assign fifo_intf_427.fifo_rd_block = 0;
    assign fifo_intf_427.fifo_wr_block = 0;
    assign fifo_intf_427.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_427;
    csv_file_dump cstatus_csv_dumper_427;
    df_fifo_monitor fifo_monitor_427;
    df_fifo_intf fifo_intf_428(clock,reset);
    assign fifo_intf_428.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_20_U.if_empty_n;
    assign fifo_intf_428.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_20_U.if_full_n;
    assign fifo_intf_428.fifo_rd_block = 0;
    assign fifo_intf_428.fifo_wr_block = 0;
    assign fifo_intf_428.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_428;
    csv_file_dump cstatus_csv_dumper_428;
    df_fifo_monitor fifo_monitor_428;
    df_fifo_intf fifo_intf_429(clock,reset);
    assign fifo_intf_429.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_20_U.if_empty_n;
    assign fifo_intf_429.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_20_U.if_full_n;
    assign fifo_intf_429.fifo_rd_block = 0;
    assign fifo_intf_429.fifo_wr_block = 0;
    assign fifo_intf_429.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_429;
    csv_file_dump cstatus_csv_dumper_429;
    df_fifo_monitor fifo_monitor_429;
    df_fifo_intf fifo_intf_430(clock,reset);
    assign fifo_intf_430.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_20_U.if_empty_n;
    assign fifo_intf_430.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_20_U.if_full_n;
    assign fifo_intf_430.fifo_rd_block = 0;
    assign fifo_intf_430.fifo_wr_block = 0;
    assign fifo_intf_430.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_430;
    csv_file_dump cstatus_csv_dumper_430;
    df_fifo_monitor fifo_monitor_430;
    df_fifo_intf fifo_intf_431(clock,reset);
    assign fifo_intf_431.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_20_U.if_empty_n;
    assign fifo_intf_431.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_20_U.if_full_n;
    assign fifo_intf_431.fifo_rd_block = 0;
    assign fifo_intf_431.fifo_wr_block = 0;
    assign fifo_intf_431.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_431;
    csv_file_dump cstatus_csv_dumper_431;
    df_fifo_monitor fifo_monitor_431;
    df_fifo_intf fifo_intf_432(clock,reset);
    assign fifo_intf_432.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_20_U.if_empty_n;
    assign fifo_intf_432.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_20_U.if_full_n;
    assign fifo_intf_432.fifo_rd_block = 0;
    assign fifo_intf_432.fifo_wr_block = 0;
    assign fifo_intf_432.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_432;
    csv_file_dump cstatus_csv_dumper_432;
    df_fifo_monitor fifo_monitor_432;
    df_fifo_intf fifo_intf_433(clock,reset);
    assign fifo_intf_433.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_20_U.if_empty_n;
    assign fifo_intf_433.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_20_U.if_full_n;
    assign fifo_intf_433.fifo_rd_block = 0;
    assign fifo_intf_433.fifo_wr_block = 0;
    assign fifo_intf_433.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_433;
    csv_file_dump cstatus_csv_dumper_433;
    df_fifo_monitor fifo_monitor_433;
    df_fifo_intf fifo_intf_434(clock,reset);
    assign fifo_intf_434.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_20_U.if_empty_n;
    assign fifo_intf_434.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_20_U.if_full_n;
    assign fifo_intf_434.fifo_rd_block = 0;
    assign fifo_intf_434.fifo_wr_block = 0;
    assign fifo_intf_434.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_434;
    csv_file_dump cstatus_csv_dumper_434;
    df_fifo_monitor fifo_monitor_434;
    df_fifo_intf fifo_intf_435(clock,reset);
    assign fifo_intf_435.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_20_U.if_empty_n;
    assign fifo_intf_435.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_20_U.if_full_n;
    assign fifo_intf_435.fifo_rd_block = 0;
    assign fifo_intf_435.fifo_wr_block = 0;
    assign fifo_intf_435.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_435;
    csv_file_dump cstatus_csv_dumper_435;
    df_fifo_monitor fifo_monitor_435;
    df_fifo_intf fifo_intf_436(clock,reset);
    assign fifo_intf_436.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_20_U.if_empty_n;
    assign fifo_intf_436.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_20_U.if_full_n;
    assign fifo_intf_436.fifo_rd_block = 0;
    assign fifo_intf_436.fifo_wr_block = 0;
    assign fifo_intf_436.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_436;
    csv_file_dump cstatus_csv_dumper_436;
    df_fifo_monitor fifo_monitor_436;
    df_fifo_intf fifo_intf_437(clock,reset);
    assign fifo_intf_437.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_20_U.if_empty_n;
    assign fifo_intf_437.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_20_U.if_full_n;
    assign fifo_intf_437.fifo_rd_block = 0;
    assign fifo_intf_437.fifo_wr_block = 0;
    assign fifo_intf_437.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_437;
    csv_file_dump cstatus_csv_dumper_437;
    df_fifo_monitor fifo_monitor_437;
    df_fifo_intf fifo_intf_438(clock,reset);
    assign fifo_intf_438.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_20_U.if_empty_n;
    assign fifo_intf_438.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_20_U.if_full_n;
    assign fifo_intf_438.fifo_rd_block = 0;
    assign fifo_intf_438.fifo_wr_block = 0;
    assign fifo_intf_438.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_438;
    csv_file_dump cstatus_csv_dumper_438;
    df_fifo_monitor fifo_monitor_438;
    df_fifo_intf fifo_intf_439(clock,reset);
    assign fifo_intf_439.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_20_U.if_empty_n;
    assign fifo_intf_439.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_20_U.if_full_n;
    assign fifo_intf_439.fifo_rd_block = 0;
    assign fifo_intf_439.fifo_wr_block = 0;
    assign fifo_intf_439.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_439;
    csv_file_dump cstatus_csv_dumper_439;
    df_fifo_monitor fifo_monitor_439;
    df_fifo_intf fifo_intf_440(clock,reset);
    assign fifo_intf_440.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_20_U.if_empty_n;
    assign fifo_intf_440.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_20_U.if_full_n;
    assign fifo_intf_440.fifo_rd_block = 0;
    assign fifo_intf_440.fifo_wr_block = 0;
    assign fifo_intf_440.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_440;
    csv_file_dump cstatus_csv_dumper_440;
    df_fifo_monitor fifo_monitor_440;
    df_fifo_intf fifo_intf_441(clock,reset);
    assign fifo_intf_441.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_20_U.if_empty_n;
    assign fifo_intf_441.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_20_U.if_full_n;
    assign fifo_intf_441.fifo_rd_block = 0;
    assign fifo_intf_441.fifo_wr_block = 0;
    assign fifo_intf_441.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_441;
    csv_file_dump cstatus_csv_dumper_441;
    df_fifo_monitor fifo_monitor_441;
    df_fifo_intf fifo_intf_442(clock,reset);
    assign fifo_intf_442.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_20_U.if_empty_n;
    assign fifo_intf_442.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_20_U.if_full_n;
    assign fifo_intf_442.fifo_rd_block = 0;
    assign fifo_intf_442.fifo_wr_block = 0;
    assign fifo_intf_442.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_442;
    csv_file_dump cstatus_csv_dumper_442;
    df_fifo_monitor fifo_monitor_442;
    df_fifo_intf fifo_intf_443(clock,reset);
    assign fifo_intf_443.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_20_U.if_empty_n;
    assign fifo_intf_443.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_20_U.if_full_n;
    assign fifo_intf_443.fifo_rd_block = 0;
    assign fifo_intf_443.fifo_wr_block = 0;
    assign fifo_intf_443.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_443;
    csv_file_dump cstatus_csv_dumper_443;
    df_fifo_monitor fifo_monitor_443;
    df_fifo_intf fifo_intf_444(clock,reset);
    assign fifo_intf_444.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_20_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_20_U.if_empty_n;
    assign fifo_intf_444.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_20_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_20_U.if_full_n;
    assign fifo_intf_444.fifo_rd_block = 0;
    assign fifo_intf_444.fifo_wr_block = 0;
    assign fifo_intf_444.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_444;
    csv_file_dump cstatus_csv_dumper_444;
    df_fifo_monitor fifo_monitor_444;
    df_fifo_intf fifo_intf_445(clock,reset);
    assign fifo_intf_445.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_21_U.if_empty_n;
    assign fifo_intf_445.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_21_U.if_full_n;
    assign fifo_intf_445.fifo_rd_block = 0;
    assign fifo_intf_445.fifo_wr_block = 0;
    assign fifo_intf_445.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_445;
    csv_file_dump cstatus_csv_dumper_445;
    df_fifo_monitor fifo_monitor_445;
    df_fifo_intf fifo_intf_446(clock,reset);
    assign fifo_intf_446.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_21_U.if_empty_n;
    assign fifo_intf_446.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_21_U.if_full_n;
    assign fifo_intf_446.fifo_rd_block = 0;
    assign fifo_intf_446.fifo_wr_block = 0;
    assign fifo_intf_446.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_446;
    csv_file_dump cstatus_csv_dumper_446;
    df_fifo_monitor fifo_monitor_446;
    df_fifo_intf fifo_intf_447(clock,reset);
    assign fifo_intf_447.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_21_U.if_empty_n;
    assign fifo_intf_447.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_21_U.if_full_n;
    assign fifo_intf_447.fifo_rd_block = 0;
    assign fifo_intf_447.fifo_wr_block = 0;
    assign fifo_intf_447.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_447;
    csv_file_dump cstatus_csv_dumper_447;
    df_fifo_monitor fifo_monitor_447;
    df_fifo_intf fifo_intf_448(clock,reset);
    assign fifo_intf_448.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_21_U.if_empty_n;
    assign fifo_intf_448.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_21_U.if_full_n;
    assign fifo_intf_448.fifo_rd_block = 0;
    assign fifo_intf_448.fifo_wr_block = 0;
    assign fifo_intf_448.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_448;
    csv_file_dump cstatus_csv_dumper_448;
    df_fifo_monitor fifo_monitor_448;
    df_fifo_intf fifo_intf_449(clock,reset);
    assign fifo_intf_449.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_21_U.if_empty_n;
    assign fifo_intf_449.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_21_U.if_full_n;
    assign fifo_intf_449.fifo_rd_block = 0;
    assign fifo_intf_449.fifo_wr_block = 0;
    assign fifo_intf_449.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_449;
    csv_file_dump cstatus_csv_dumper_449;
    df_fifo_monitor fifo_monitor_449;
    df_fifo_intf fifo_intf_450(clock,reset);
    assign fifo_intf_450.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_21_U.if_empty_n;
    assign fifo_intf_450.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_21_U.if_full_n;
    assign fifo_intf_450.fifo_rd_block = 0;
    assign fifo_intf_450.fifo_wr_block = 0;
    assign fifo_intf_450.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_450;
    csv_file_dump cstatus_csv_dumper_450;
    df_fifo_monitor fifo_monitor_450;
    df_fifo_intf fifo_intf_451(clock,reset);
    assign fifo_intf_451.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_21_U.if_empty_n;
    assign fifo_intf_451.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_21_U.if_full_n;
    assign fifo_intf_451.fifo_rd_block = 0;
    assign fifo_intf_451.fifo_wr_block = 0;
    assign fifo_intf_451.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_451;
    csv_file_dump cstatus_csv_dumper_451;
    df_fifo_monitor fifo_monitor_451;
    df_fifo_intf fifo_intf_452(clock,reset);
    assign fifo_intf_452.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_21_U.if_empty_n;
    assign fifo_intf_452.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_21_U.if_full_n;
    assign fifo_intf_452.fifo_rd_block = 0;
    assign fifo_intf_452.fifo_wr_block = 0;
    assign fifo_intf_452.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_452;
    csv_file_dump cstatus_csv_dumper_452;
    df_fifo_monitor fifo_monitor_452;
    df_fifo_intf fifo_intf_453(clock,reset);
    assign fifo_intf_453.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_21_U.if_empty_n;
    assign fifo_intf_453.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_21_U.if_full_n;
    assign fifo_intf_453.fifo_rd_block = 0;
    assign fifo_intf_453.fifo_wr_block = 0;
    assign fifo_intf_453.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_453;
    csv_file_dump cstatus_csv_dumper_453;
    df_fifo_monitor fifo_monitor_453;
    df_fifo_intf fifo_intf_454(clock,reset);
    assign fifo_intf_454.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_21_U.if_empty_n;
    assign fifo_intf_454.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_21_U.if_full_n;
    assign fifo_intf_454.fifo_rd_block = 0;
    assign fifo_intf_454.fifo_wr_block = 0;
    assign fifo_intf_454.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_454;
    csv_file_dump cstatus_csv_dumper_454;
    df_fifo_monitor fifo_monitor_454;
    df_fifo_intf fifo_intf_455(clock,reset);
    assign fifo_intf_455.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_21_U.if_empty_n;
    assign fifo_intf_455.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_21_U.if_full_n;
    assign fifo_intf_455.fifo_rd_block = 0;
    assign fifo_intf_455.fifo_wr_block = 0;
    assign fifo_intf_455.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_455;
    csv_file_dump cstatus_csv_dumper_455;
    df_fifo_monitor fifo_monitor_455;
    df_fifo_intf fifo_intf_456(clock,reset);
    assign fifo_intf_456.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_21_U.if_empty_n;
    assign fifo_intf_456.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_21_U.if_full_n;
    assign fifo_intf_456.fifo_rd_block = 0;
    assign fifo_intf_456.fifo_wr_block = 0;
    assign fifo_intf_456.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_456;
    csv_file_dump cstatus_csv_dumper_456;
    df_fifo_monitor fifo_monitor_456;
    df_fifo_intf fifo_intf_457(clock,reset);
    assign fifo_intf_457.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_21_U.if_empty_n;
    assign fifo_intf_457.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_21_U.if_full_n;
    assign fifo_intf_457.fifo_rd_block = 0;
    assign fifo_intf_457.fifo_wr_block = 0;
    assign fifo_intf_457.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_457;
    csv_file_dump cstatus_csv_dumper_457;
    df_fifo_monitor fifo_monitor_457;
    df_fifo_intf fifo_intf_458(clock,reset);
    assign fifo_intf_458.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_21_U.if_empty_n;
    assign fifo_intf_458.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_21_U.if_full_n;
    assign fifo_intf_458.fifo_rd_block = 0;
    assign fifo_intf_458.fifo_wr_block = 0;
    assign fifo_intf_458.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_458;
    csv_file_dump cstatus_csv_dumper_458;
    df_fifo_monitor fifo_monitor_458;
    df_fifo_intf fifo_intf_459(clock,reset);
    assign fifo_intf_459.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_21_U.if_empty_n;
    assign fifo_intf_459.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_21_U.if_full_n;
    assign fifo_intf_459.fifo_rd_block = 0;
    assign fifo_intf_459.fifo_wr_block = 0;
    assign fifo_intf_459.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_459;
    csv_file_dump cstatus_csv_dumper_459;
    df_fifo_monitor fifo_monitor_459;
    df_fifo_intf fifo_intf_460(clock,reset);
    assign fifo_intf_460.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_21_U.if_empty_n;
    assign fifo_intf_460.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_21_U.if_full_n;
    assign fifo_intf_460.fifo_rd_block = 0;
    assign fifo_intf_460.fifo_wr_block = 0;
    assign fifo_intf_460.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_460;
    csv_file_dump cstatus_csv_dumper_460;
    df_fifo_monitor fifo_monitor_460;
    df_fifo_intf fifo_intf_461(clock,reset);
    assign fifo_intf_461.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_21_U.if_empty_n;
    assign fifo_intf_461.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_21_U.if_full_n;
    assign fifo_intf_461.fifo_rd_block = 0;
    assign fifo_intf_461.fifo_wr_block = 0;
    assign fifo_intf_461.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_461;
    csv_file_dump cstatus_csv_dumper_461;
    df_fifo_monitor fifo_monitor_461;
    df_fifo_intf fifo_intf_462(clock,reset);
    assign fifo_intf_462.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_21_U.if_empty_n;
    assign fifo_intf_462.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_21_U.if_full_n;
    assign fifo_intf_462.fifo_rd_block = 0;
    assign fifo_intf_462.fifo_wr_block = 0;
    assign fifo_intf_462.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_462;
    csv_file_dump cstatus_csv_dumper_462;
    df_fifo_monitor fifo_monitor_462;
    df_fifo_intf fifo_intf_463(clock,reset);
    assign fifo_intf_463.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_21_U.if_empty_n;
    assign fifo_intf_463.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_21_U.if_full_n;
    assign fifo_intf_463.fifo_rd_block = 0;
    assign fifo_intf_463.fifo_wr_block = 0;
    assign fifo_intf_463.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_463;
    csv_file_dump cstatus_csv_dumper_463;
    df_fifo_monitor fifo_monitor_463;
    df_fifo_intf fifo_intf_464(clock,reset);
    assign fifo_intf_464.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_21_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_21_U.if_empty_n;
    assign fifo_intf_464.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_21_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_21_U.if_full_n;
    assign fifo_intf_464.fifo_rd_block = 0;
    assign fifo_intf_464.fifo_wr_block = 0;
    assign fifo_intf_464.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_464;
    csv_file_dump cstatus_csv_dumper_464;
    df_fifo_monitor fifo_monitor_464;
    df_fifo_intf fifo_intf_465(clock,reset);
    assign fifo_intf_465.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_22_U.if_empty_n;
    assign fifo_intf_465.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_22_U.if_full_n;
    assign fifo_intf_465.fifo_rd_block = 0;
    assign fifo_intf_465.fifo_wr_block = 0;
    assign fifo_intf_465.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_465;
    csv_file_dump cstatus_csv_dumper_465;
    df_fifo_monitor fifo_monitor_465;
    df_fifo_intf fifo_intf_466(clock,reset);
    assign fifo_intf_466.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_22_U.if_empty_n;
    assign fifo_intf_466.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_22_U.if_full_n;
    assign fifo_intf_466.fifo_rd_block = 0;
    assign fifo_intf_466.fifo_wr_block = 0;
    assign fifo_intf_466.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_466;
    csv_file_dump cstatus_csv_dumper_466;
    df_fifo_monitor fifo_monitor_466;
    df_fifo_intf fifo_intf_467(clock,reset);
    assign fifo_intf_467.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_22_U.if_empty_n;
    assign fifo_intf_467.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_22_U.if_full_n;
    assign fifo_intf_467.fifo_rd_block = 0;
    assign fifo_intf_467.fifo_wr_block = 0;
    assign fifo_intf_467.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_467;
    csv_file_dump cstatus_csv_dumper_467;
    df_fifo_monitor fifo_monitor_467;
    df_fifo_intf fifo_intf_468(clock,reset);
    assign fifo_intf_468.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_22_U.if_empty_n;
    assign fifo_intf_468.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_22_U.if_full_n;
    assign fifo_intf_468.fifo_rd_block = 0;
    assign fifo_intf_468.fifo_wr_block = 0;
    assign fifo_intf_468.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_468;
    csv_file_dump cstatus_csv_dumper_468;
    df_fifo_monitor fifo_monitor_468;
    df_fifo_intf fifo_intf_469(clock,reset);
    assign fifo_intf_469.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_22_U.if_empty_n;
    assign fifo_intf_469.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_22_U.if_full_n;
    assign fifo_intf_469.fifo_rd_block = 0;
    assign fifo_intf_469.fifo_wr_block = 0;
    assign fifo_intf_469.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_469;
    csv_file_dump cstatus_csv_dumper_469;
    df_fifo_monitor fifo_monitor_469;
    df_fifo_intf fifo_intf_470(clock,reset);
    assign fifo_intf_470.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_22_U.if_empty_n;
    assign fifo_intf_470.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_22_U.if_full_n;
    assign fifo_intf_470.fifo_rd_block = 0;
    assign fifo_intf_470.fifo_wr_block = 0;
    assign fifo_intf_470.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_470;
    csv_file_dump cstatus_csv_dumper_470;
    df_fifo_monitor fifo_monitor_470;
    df_fifo_intf fifo_intf_471(clock,reset);
    assign fifo_intf_471.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_22_U.if_empty_n;
    assign fifo_intf_471.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_22_U.if_full_n;
    assign fifo_intf_471.fifo_rd_block = 0;
    assign fifo_intf_471.fifo_wr_block = 0;
    assign fifo_intf_471.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_471;
    csv_file_dump cstatus_csv_dumper_471;
    df_fifo_monitor fifo_monitor_471;
    df_fifo_intf fifo_intf_472(clock,reset);
    assign fifo_intf_472.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_22_U.if_empty_n;
    assign fifo_intf_472.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_22_U.if_full_n;
    assign fifo_intf_472.fifo_rd_block = 0;
    assign fifo_intf_472.fifo_wr_block = 0;
    assign fifo_intf_472.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_472;
    csv_file_dump cstatus_csv_dumper_472;
    df_fifo_monitor fifo_monitor_472;
    df_fifo_intf fifo_intf_473(clock,reset);
    assign fifo_intf_473.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_22_U.if_empty_n;
    assign fifo_intf_473.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_22_U.if_full_n;
    assign fifo_intf_473.fifo_rd_block = 0;
    assign fifo_intf_473.fifo_wr_block = 0;
    assign fifo_intf_473.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_473;
    csv_file_dump cstatus_csv_dumper_473;
    df_fifo_monitor fifo_monitor_473;
    df_fifo_intf fifo_intf_474(clock,reset);
    assign fifo_intf_474.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_22_U.if_empty_n;
    assign fifo_intf_474.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_22_U.if_full_n;
    assign fifo_intf_474.fifo_rd_block = 0;
    assign fifo_intf_474.fifo_wr_block = 0;
    assign fifo_intf_474.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_474;
    csv_file_dump cstatus_csv_dumper_474;
    df_fifo_monitor fifo_monitor_474;
    df_fifo_intf fifo_intf_475(clock,reset);
    assign fifo_intf_475.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_22_U.if_empty_n;
    assign fifo_intf_475.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_22_U.if_full_n;
    assign fifo_intf_475.fifo_rd_block = 0;
    assign fifo_intf_475.fifo_wr_block = 0;
    assign fifo_intf_475.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_475;
    csv_file_dump cstatus_csv_dumper_475;
    df_fifo_monitor fifo_monitor_475;
    df_fifo_intf fifo_intf_476(clock,reset);
    assign fifo_intf_476.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_22_U.if_empty_n;
    assign fifo_intf_476.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_22_U.if_full_n;
    assign fifo_intf_476.fifo_rd_block = 0;
    assign fifo_intf_476.fifo_wr_block = 0;
    assign fifo_intf_476.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_476;
    csv_file_dump cstatus_csv_dumper_476;
    df_fifo_monitor fifo_monitor_476;
    df_fifo_intf fifo_intf_477(clock,reset);
    assign fifo_intf_477.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_22_U.if_empty_n;
    assign fifo_intf_477.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_22_U.if_full_n;
    assign fifo_intf_477.fifo_rd_block = 0;
    assign fifo_intf_477.fifo_wr_block = 0;
    assign fifo_intf_477.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_477;
    csv_file_dump cstatus_csv_dumper_477;
    df_fifo_monitor fifo_monitor_477;
    df_fifo_intf fifo_intf_478(clock,reset);
    assign fifo_intf_478.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_22_U.if_empty_n;
    assign fifo_intf_478.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_22_U.if_full_n;
    assign fifo_intf_478.fifo_rd_block = 0;
    assign fifo_intf_478.fifo_wr_block = 0;
    assign fifo_intf_478.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_478;
    csv_file_dump cstatus_csv_dumper_478;
    df_fifo_monitor fifo_monitor_478;
    df_fifo_intf fifo_intf_479(clock,reset);
    assign fifo_intf_479.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_22_U.if_empty_n;
    assign fifo_intf_479.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_22_U.if_full_n;
    assign fifo_intf_479.fifo_rd_block = 0;
    assign fifo_intf_479.fifo_wr_block = 0;
    assign fifo_intf_479.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_479;
    csv_file_dump cstatus_csv_dumper_479;
    df_fifo_monitor fifo_monitor_479;
    df_fifo_intf fifo_intf_480(clock,reset);
    assign fifo_intf_480.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_22_U.if_empty_n;
    assign fifo_intf_480.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_22_U.if_full_n;
    assign fifo_intf_480.fifo_rd_block = 0;
    assign fifo_intf_480.fifo_wr_block = 0;
    assign fifo_intf_480.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_480;
    csv_file_dump cstatus_csv_dumper_480;
    df_fifo_monitor fifo_monitor_480;
    df_fifo_intf fifo_intf_481(clock,reset);
    assign fifo_intf_481.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_22_U.if_empty_n;
    assign fifo_intf_481.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_22_U.if_full_n;
    assign fifo_intf_481.fifo_rd_block = 0;
    assign fifo_intf_481.fifo_wr_block = 0;
    assign fifo_intf_481.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_481;
    csv_file_dump cstatus_csv_dumper_481;
    df_fifo_monitor fifo_monitor_481;
    df_fifo_intf fifo_intf_482(clock,reset);
    assign fifo_intf_482.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_22_U.if_empty_n;
    assign fifo_intf_482.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_22_U.if_full_n;
    assign fifo_intf_482.fifo_rd_block = 0;
    assign fifo_intf_482.fifo_wr_block = 0;
    assign fifo_intf_482.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_482;
    csv_file_dump cstatus_csv_dumper_482;
    df_fifo_monitor fifo_monitor_482;
    df_fifo_intf fifo_intf_483(clock,reset);
    assign fifo_intf_483.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_22_U.if_empty_n;
    assign fifo_intf_483.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_22_U.if_full_n;
    assign fifo_intf_483.fifo_rd_block = 0;
    assign fifo_intf_483.fifo_wr_block = 0;
    assign fifo_intf_483.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_483;
    csv_file_dump cstatus_csv_dumper_483;
    df_fifo_monitor fifo_monitor_483;
    df_fifo_intf fifo_intf_484(clock,reset);
    assign fifo_intf_484.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_22_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_22_U.if_empty_n;
    assign fifo_intf_484.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_22_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_22_U.if_full_n;
    assign fifo_intf_484.fifo_rd_block = 0;
    assign fifo_intf_484.fifo_wr_block = 0;
    assign fifo_intf_484.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_484;
    csv_file_dump cstatus_csv_dumper_484;
    df_fifo_monitor fifo_monitor_484;
    df_fifo_intf fifo_intf_485(clock,reset);
    assign fifo_intf_485.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_23_U.if_empty_n;
    assign fifo_intf_485.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_23_U.if_full_n;
    assign fifo_intf_485.fifo_rd_block = 0;
    assign fifo_intf_485.fifo_wr_block = 0;
    assign fifo_intf_485.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_485;
    csv_file_dump cstatus_csv_dumper_485;
    df_fifo_monitor fifo_monitor_485;
    df_fifo_intf fifo_intf_486(clock,reset);
    assign fifo_intf_486.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_23_U.if_empty_n;
    assign fifo_intf_486.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_23_U.if_full_n;
    assign fifo_intf_486.fifo_rd_block = 0;
    assign fifo_intf_486.fifo_wr_block = 0;
    assign fifo_intf_486.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_486;
    csv_file_dump cstatus_csv_dumper_486;
    df_fifo_monitor fifo_monitor_486;
    df_fifo_intf fifo_intf_487(clock,reset);
    assign fifo_intf_487.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_23_U.if_empty_n;
    assign fifo_intf_487.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_23_U.if_full_n;
    assign fifo_intf_487.fifo_rd_block = 0;
    assign fifo_intf_487.fifo_wr_block = 0;
    assign fifo_intf_487.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_487;
    csv_file_dump cstatus_csv_dumper_487;
    df_fifo_monitor fifo_monitor_487;
    df_fifo_intf fifo_intf_488(clock,reset);
    assign fifo_intf_488.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_23_U.if_empty_n;
    assign fifo_intf_488.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_23_U.if_full_n;
    assign fifo_intf_488.fifo_rd_block = 0;
    assign fifo_intf_488.fifo_wr_block = 0;
    assign fifo_intf_488.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_488;
    csv_file_dump cstatus_csv_dumper_488;
    df_fifo_monitor fifo_monitor_488;
    df_fifo_intf fifo_intf_489(clock,reset);
    assign fifo_intf_489.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_23_U.if_empty_n;
    assign fifo_intf_489.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_23_U.if_full_n;
    assign fifo_intf_489.fifo_rd_block = 0;
    assign fifo_intf_489.fifo_wr_block = 0;
    assign fifo_intf_489.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_489;
    csv_file_dump cstatus_csv_dumper_489;
    df_fifo_monitor fifo_monitor_489;
    df_fifo_intf fifo_intf_490(clock,reset);
    assign fifo_intf_490.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_23_U.if_empty_n;
    assign fifo_intf_490.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_23_U.if_full_n;
    assign fifo_intf_490.fifo_rd_block = 0;
    assign fifo_intf_490.fifo_wr_block = 0;
    assign fifo_intf_490.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_490;
    csv_file_dump cstatus_csv_dumper_490;
    df_fifo_monitor fifo_monitor_490;
    df_fifo_intf fifo_intf_491(clock,reset);
    assign fifo_intf_491.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_23_U.if_empty_n;
    assign fifo_intf_491.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_23_U.if_full_n;
    assign fifo_intf_491.fifo_rd_block = 0;
    assign fifo_intf_491.fifo_wr_block = 0;
    assign fifo_intf_491.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_491;
    csv_file_dump cstatus_csv_dumper_491;
    df_fifo_monitor fifo_monitor_491;
    df_fifo_intf fifo_intf_492(clock,reset);
    assign fifo_intf_492.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_23_U.if_empty_n;
    assign fifo_intf_492.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_23_U.if_full_n;
    assign fifo_intf_492.fifo_rd_block = 0;
    assign fifo_intf_492.fifo_wr_block = 0;
    assign fifo_intf_492.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_492;
    csv_file_dump cstatus_csv_dumper_492;
    df_fifo_monitor fifo_monitor_492;
    df_fifo_intf fifo_intf_493(clock,reset);
    assign fifo_intf_493.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_23_U.if_empty_n;
    assign fifo_intf_493.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_23_U.if_full_n;
    assign fifo_intf_493.fifo_rd_block = 0;
    assign fifo_intf_493.fifo_wr_block = 0;
    assign fifo_intf_493.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_493;
    csv_file_dump cstatus_csv_dumper_493;
    df_fifo_monitor fifo_monitor_493;
    df_fifo_intf fifo_intf_494(clock,reset);
    assign fifo_intf_494.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_23_U.if_empty_n;
    assign fifo_intf_494.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_23_U.if_full_n;
    assign fifo_intf_494.fifo_rd_block = 0;
    assign fifo_intf_494.fifo_wr_block = 0;
    assign fifo_intf_494.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_494;
    csv_file_dump cstatus_csv_dumper_494;
    df_fifo_monitor fifo_monitor_494;
    df_fifo_intf fifo_intf_495(clock,reset);
    assign fifo_intf_495.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_23_U.if_empty_n;
    assign fifo_intf_495.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_23_U.if_full_n;
    assign fifo_intf_495.fifo_rd_block = 0;
    assign fifo_intf_495.fifo_wr_block = 0;
    assign fifo_intf_495.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_495;
    csv_file_dump cstatus_csv_dumper_495;
    df_fifo_monitor fifo_monitor_495;
    df_fifo_intf fifo_intf_496(clock,reset);
    assign fifo_intf_496.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_23_U.if_empty_n;
    assign fifo_intf_496.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_23_U.if_full_n;
    assign fifo_intf_496.fifo_rd_block = 0;
    assign fifo_intf_496.fifo_wr_block = 0;
    assign fifo_intf_496.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_496;
    csv_file_dump cstatus_csv_dumper_496;
    df_fifo_monitor fifo_monitor_496;
    df_fifo_intf fifo_intf_497(clock,reset);
    assign fifo_intf_497.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_23_U.if_empty_n;
    assign fifo_intf_497.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_23_U.if_full_n;
    assign fifo_intf_497.fifo_rd_block = 0;
    assign fifo_intf_497.fifo_wr_block = 0;
    assign fifo_intf_497.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_497;
    csv_file_dump cstatus_csv_dumper_497;
    df_fifo_monitor fifo_monitor_497;
    df_fifo_intf fifo_intf_498(clock,reset);
    assign fifo_intf_498.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_23_U.if_empty_n;
    assign fifo_intf_498.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_23_U.if_full_n;
    assign fifo_intf_498.fifo_rd_block = 0;
    assign fifo_intf_498.fifo_wr_block = 0;
    assign fifo_intf_498.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_498;
    csv_file_dump cstatus_csv_dumper_498;
    df_fifo_monitor fifo_monitor_498;
    df_fifo_intf fifo_intf_499(clock,reset);
    assign fifo_intf_499.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_23_U.if_empty_n;
    assign fifo_intf_499.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_23_U.if_full_n;
    assign fifo_intf_499.fifo_rd_block = 0;
    assign fifo_intf_499.fifo_wr_block = 0;
    assign fifo_intf_499.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_499;
    csv_file_dump cstatus_csv_dumper_499;
    df_fifo_monitor fifo_monitor_499;
    df_fifo_intf fifo_intf_500(clock,reset);
    assign fifo_intf_500.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_23_U.if_empty_n;
    assign fifo_intf_500.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_23_U.if_full_n;
    assign fifo_intf_500.fifo_rd_block = 0;
    assign fifo_intf_500.fifo_wr_block = 0;
    assign fifo_intf_500.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_500;
    csv_file_dump cstatus_csv_dumper_500;
    df_fifo_monitor fifo_monitor_500;
    df_fifo_intf fifo_intf_501(clock,reset);
    assign fifo_intf_501.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_23_U.if_empty_n;
    assign fifo_intf_501.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_23_U.if_full_n;
    assign fifo_intf_501.fifo_rd_block = 0;
    assign fifo_intf_501.fifo_wr_block = 0;
    assign fifo_intf_501.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_501;
    csv_file_dump cstatus_csv_dumper_501;
    df_fifo_monitor fifo_monitor_501;
    df_fifo_intf fifo_intf_502(clock,reset);
    assign fifo_intf_502.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_23_U.if_empty_n;
    assign fifo_intf_502.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_23_U.if_full_n;
    assign fifo_intf_502.fifo_rd_block = 0;
    assign fifo_intf_502.fifo_wr_block = 0;
    assign fifo_intf_502.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_502;
    csv_file_dump cstatus_csv_dumper_502;
    df_fifo_monitor fifo_monitor_502;
    df_fifo_intf fifo_intf_503(clock,reset);
    assign fifo_intf_503.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_23_U.if_empty_n;
    assign fifo_intf_503.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_23_U.if_full_n;
    assign fifo_intf_503.fifo_rd_block = 0;
    assign fifo_intf_503.fifo_wr_block = 0;
    assign fifo_intf_503.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_503;
    csv_file_dump cstatus_csv_dumper_503;
    df_fifo_monitor fifo_monitor_503;
    df_fifo_intf fifo_intf_504(clock,reset);
    assign fifo_intf_504.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_23_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_23_U.if_empty_n;
    assign fifo_intf_504.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_23_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_23_U.if_full_n;
    assign fifo_intf_504.fifo_rd_block = 0;
    assign fifo_intf_504.fifo_wr_block = 0;
    assign fifo_intf_504.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_504;
    csv_file_dump cstatus_csv_dumper_504;
    df_fifo_monitor fifo_monitor_504;
    df_fifo_intf fifo_intf_505(clock,reset);
    assign fifo_intf_505.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_24_U.if_empty_n;
    assign fifo_intf_505.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_24_U.if_full_n;
    assign fifo_intf_505.fifo_rd_block = 0;
    assign fifo_intf_505.fifo_wr_block = 0;
    assign fifo_intf_505.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_505;
    csv_file_dump cstatus_csv_dumper_505;
    df_fifo_monitor fifo_monitor_505;
    df_fifo_intf fifo_intf_506(clock,reset);
    assign fifo_intf_506.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_24_U.if_empty_n;
    assign fifo_intf_506.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_24_U.if_full_n;
    assign fifo_intf_506.fifo_rd_block = 0;
    assign fifo_intf_506.fifo_wr_block = 0;
    assign fifo_intf_506.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_506;
    csv_file_dump cstatus_csv_dumper_506;
    df_fifo_monitor fifo_monitor_506;
    df_fifo_intf fifo_intf_507(clock,reset);
    assign fifo_intf_507.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_24_U.if_empty_n;
    assign fifo_intf_507.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_24_U.if_full_n;
    assign fifo_intf_507.fifo_rd_block = 0;
    assign fifo_intf_507.fifo_wr_block = 0;
    assign fifo_intf_507.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_507;
    csv_file_dump cstatus_csv_dumper_507;
    df_fifo_monitor fifo_monitor_507;
    df_fifo_intf fifo_intf_508(clock,reset);
    assign fifo_intf_508.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_24_U.if_empty_n;
    assign fifo_intf_508.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_24_U.if_full_n;
    assign fifo_intf_508.fifo_rd_block = 0;
    assign fifo_intf_508.fifo_wr_block = 0;
    assign fifo_intf_508.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_508;
    csv_file_dump cstatus_csv_dumper_508;
    df_fifo_monitor fifo_monitor_508;
    df_fifo_intf fifo_intf_509(clock,reset);
    assign fifo_intf_509.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_24_U.if_empty_n;
    assign fifo_intf_509.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_24_U.if_full_n;
    assign fifo_intf_509.fifo_rd_block = 0;
    assign fifo_intf_509.fifo_wr_block = 0;
    assign fifo_intf_509.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_509;
    csv_file_dump cstatus_csv_dumper_509;
    df_fifo_monitor fifo_monitor_509;
    df_fifo_intf fifo_intf_510(clock,reset);
    assign fifo_intf_510.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_24_U.if_empty_n;
    assign fifo_intf_510.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_24_U.if_full_n;
    assign fifo_intf_510.fifo_rd_block = 0;
    assign fifo_intf_510.fifo_wr_block = 0;
    assign fifo_intf_510.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_510;
    csv_file_dump cstatus_csv_dumper_510;
    df_fifo_monitor fifo_monitor_510;
    df_fifo_intf fifo_intf_511(clock,reset);
    assign fifo_intf_511.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_24_U.if_empty_n;
    assign fifo_intf_511.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_24_U.if_full_n;
    assign fifo_intf_511.fifo_rd_block = 0;
    assign fifo_intf_511.fifo_wr_block = 0;
    assign fifo_intf_511.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_511;
    csv_file_dump cstatus_csv_dumper_511;
    df_fifo_monitor fifo_monitor_511;
    df_fifo_intf fifo_intf_512(clock,reset);
    assign fifo_intf_512.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_24_U.if_empty_n;
    assign fifo_intf_512.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_24_U.if_full_n;
    assign fifo_intf_512.fifo_rd_block = 0;
    assign fifo_intf_512.fifo_wr_block = 0;
    assign fifo_intf_512.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_512;
    csv_file_dump cstatus_csv_dumper_512;
    df_fifo_monitor fifo_monitor_512;
    df_fifo_intf fifo_intf_513(clock,reset);
    assign fifo_intf_513.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_24_U.if_empty_n;
    assign fifo_intf_513.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_24_U.if_full_n;
    assign fifo_intf_513.fifo_rd_block = 0;
    assign fifo_intf_513.fifo_wr_block = 0;
    assign fifo_intf_513.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_513;
    csv_file_dump cstatus_csv_dumper_513;
    df_fifo_monitor fifo_monitor_513;
    df_fifo_intf fifo_intf_514(clock,reset);
    assign fifo_intf_514.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_24_U.if_empty_n;
    assign fifo_intf_514.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_24_U.if_full_n;
    assign fifo_intf_514.fifo_rd_block = 0;
    assign fifo_intf_514.fifo_wr_block = 0;
    assign fifo_intf_514.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_514;
    csv_file_dump cstatus_csv_dumper_514;
    df_fifo_monitor fifo_monitor_514;
    df_fifo_intf fifo_intf_515(clock,reset);
    assign fifo_intf_515.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_24_U.if_empty_n;
    assign fifo_intf_515.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_24_U.if_full_n;
    assign fifo_intf_515.fifo_rd_block = 0;
    assign fifo_intf_515.fifo_wr_block = 0;
    assign fifo_intf_515.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_515;
    csv_file_dump cstatus_csv_dumper_515;
    df_fifo_monitor fifo_monitor_515;
    df_fifo_intf fifo_intf_516(clock,reset);
    assign fifo_intf_516.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_24_U.if_empty_n;
    assign fifo_intf_516.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_24_U.if_full_n;
    assign fifo_intf_516.fifo_rd_block = 0;
    assign fifo_intf_516.fifo_wr_block = 0;
    assign fifo_intf_516.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_516;
    csv_file_dump cstatus_csv_dumper_516;
    df_fifo_monitor fifo_monitor_516;
    df_fifo_intf fifo_intf_517(clock,reset);
    assign fifo_intf_517.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_24_U.if_empty_n;
    assign fifo_intf_517.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_24_U.if_full_n;
    assign fifo_intf_517.fifo_rd_block = 0;
    assign fifo_intf_517.fifo_wr_block = 0;
    assign fifo_intf_517.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_517;
    csv_file_dump cstatus_csv_dumper_517;
    df_fifo_monitor fifo_monitor_517;
    df_fifo_intf fifo_intf_518(clock,reset);
    assign fifo_intf_518.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_24_U.if_empty_n;
    assign fifo_intf_518.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_24_U.if_full_n;
    assign fifo_intf_518.fifo_rd_block = 0;
    assign fifo_intf_518.fifo_wr_block = 0;
    assign fifo_intf_518.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_518;
    csv_file_dump cstatus_csv_dumper_518;
    df_fifo_monitor fifo_monitor_518;
    df_fifo_intf fifo_intf_519(clock,reset);
    assign fifo_intf_519.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_24_U.if_empty_n;
    assign fifo_intf_519.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_24_U.if_full_n;
    assign fifo_intf_519.fifo_rd_block = 0;
    assign fifo_intf_519.fifo_wr_block = 0;
    assign fifo_intf_519.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_519;
    csv_file_dump cstatus_csv_dumper_519;
    df_fifo_monitor fifo_monitor_519;
    df_fifo_intf fifo_intf_520(clock,reset);
    assign fifo_intf_520.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_24_U.if_empty_n;
    assign fifo_intf_520.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_24_U.if_full_n;
    assign fifo_intf_520.fifo_rd_block = 0;
    assign fifo_intf_520.fifo_wr_block = 0;
    assign fifo_intf_520.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_520;
    csv_file_dump cstatus_csv_dumper_520;
    df_fifo_monitor fifo_monitor_520;
    df_fifo_intf fifo_intf_521(clock,reset);
    assign fifo_intf_521.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_24_U.if_empty_n;
    assign fifo_intf_521.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_24_U.if_full_n;
    assign fifo_intf_521.fifo_rd_block = 0;
    assign fifo_intf_521.fifo_wr_block = 0;
    assign fifo_intf_521.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_521;
    csv_file_dump cstatus_csv_dumper_521;
    df_fifo_monitor fifo_monitor_521;
    df_fifo_intf fifo_intf_522(clock,reset);
    assign fifo_intf_522.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_24_U.if_empty_n;
    assign fifo_intf_522.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_24_U.if_full_n;
    assign fifo_intf_522.fifo_rd_block = 0;
    assign fifo_intf_522.fifo_wr_block = 0;
    assign fifo_intf_522.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_522;
    csv_file_dump cstatus_csv_dumper_522;
    df_fifo_monitor fifo_monitor_522;
    df_fifo_intf fifo_intf_523(clock,reset);
    assign fifo_intf_523.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_24_U.if_empty_n;
    assign fifo_intf_523.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_24_U.if_full_n;
    assign fifo_intf_523.fifo_rd_block = 0;
    assign fifo_intf_523.fifo_wr_block = 0;
    assign fifo_intf_523.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_523;
    csv_file_dump cstatus_csv_dumper_523;
    df_fifo_monitor fifo_monitor_523;
    df_fifo_intf fifo_intf_524(clock,reset);
    assign fifo_intf_524.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_24_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_24_U.if_empty_n;
    assign fifo_intf_524.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_24_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_24_U.if_full_n;
    assign fifo_intf_524.fifo_rd_block = 0;
    assign fifo_intf_524.fifo_wr_block = 0;
    assign fifo_intf_524.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_524;
    csv_file_dump cstatus_csv_dumper_524;
    df_fifo_monitor fifo_monitor_524;
    df_fifo_intf fifo_intf_525(clock,reset);
    assign fifo_intf_525.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_25_U.if_empty_n;
    assign fifo_intf_525.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_25_U.if_full_n;
    assign fifo_intf_525.fifo_rd_block = 0;
    assign fifo_intf_525.fifo_wr_block = 0;
    assign fifo_intf_525.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_525;
    csv_file_dump cstatus_csv_dumper_525;
    df_fifo_monitor fifo_monitor_525;
    df_fifo_intf fifo_intf_526(clock,reset);
    assign fifo_intf_526.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_25_U.if_empty_n;
    assign fifo_intf_526.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_25_U.if_full_n;
    assign fifo_intf_526.fifo_rd_block = 0;
    assign fifo_intf_526.fifo_wr_block = 0;
    assign fifo_intf_526.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_526;
    csv_file_dump cstatus_csv_dumper_526;
    df_fifo_monitor fifo_monitor_526;
    df_fifo_intf fifo_intf_527(clock,reset);
    assign fifo_intf_527.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_25_U.if_empty_n;
    assign fifo_intf_527.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_25_U.if_full_n;
    assign fifo_intf_527.fifo_rd_block = 0;
    assign fifo_intf_527.fifo_wr_block = 0;
    assign fifo_intf_527.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_527;
    csv_file_dump cstatus_csv_dumper_527;
    df_fifo_monitor fifo_monitor_527;
    df_fifo_intf fifo_intf_528(clock,reset);
    assign fifo_intf_528.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_25_U.if_empty_n;
    assign fifo_intf_528.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_25_U.if_full_n;
    assign fifo_intf_528.fifo_rd_block = 0;
    assign fifo_intf_528.fifo_wr_block = 0;
    assign fifo_intf_528.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_528;
    csv_file_dump cstatus_csv_dumper_528;
    df_fifo_monitor fifo_monitor_528;
    df_fifo_intf fifo_intf_529(clock,reset);
    assign fifo_intf_529.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_25_U.if_empty_n;
    assign fifo_intf_529.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_25_U.if_full_n;
    assign fifo_intf_529.fifo_rd_block = 0;
    assign fifo_intf_529.fifo_wr_block = 0;
    assign fifo_intf_529.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_529;
    csv_file_dump cstatus_csv_dumper_529;
    df_fifo_monitor fifo_monitor_529;
    df_fifo_intf fifo_intf_530(clock,reset);
    assign fifo_intf_530.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_25_U.if_empty_n;
    assign fifo_intf_530.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_25_U.if_full_n;
    assign fifo_intf_530.fifo_rd_block = 0;
    assign fifo_intf_530.fifo_wr_block = 0;
    assign fifo_intf_530.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_530;
    csv_file_dump cstatus_csv_dumper_530;
    df_fifo_monitor fifo_monitor_530;
    df_fifo_intf fifo_intf_531(clock,reset);
    assign fifo_intf_531.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_25_U.if_empty_n;
    assign fifo_intf_531.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_25_U.if_full_n;
    assign fifo_intf_531.fifo_rd_block = 0;
    assign fifo_intf_531.fifo_wr_block = 0;
    assign fifo_intf_531.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_531;
    csv_file_dump cstatus_csv_dumper_531;
    df_fifo_monitor fifo_monitor_531;
    df_fifo_intf fifo_intf_532(clock,reset);
    assign fifo_intf_532.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_25_U.if_empty_n;
    assign fifo_intf_532.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_25_U.if_full_n;
    assign fifo_intf_532.fifo_rd_block = 0;
    assign fifo_intf_532.fifo_wr_block = 0;
    assign fifo_intf_532.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_532;
    csv_file_dump cstatus_csv_dumper_532;
    df_fifo_monitor fifo_monitor_532;
    df_fifo_intf fifo_intf_533(clock,reset);
    assign fifo_intf_533.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_25_U.if_empty_n;
    assign fifo_intf_533.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_25_U.if_full_n;
    assign fifo_intf_533.fifo_rd_block = 0;
    assign fifo_intf_533.fifo_wr_block = 0;
    assign fifo_intf_533.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_533;
    csv_file_dump cstatus_csv_dumper_533;
    df_fifo_monitor fifo_monitor_533;
    df_fifo_intf fifo_intf_534(clock,reset);
    assign fifo_intf_534.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_25_U.if_empty_n;
    assign fifo_intf_534.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_25_U.if_full_n;
    assign fifo_intf_534.fifo_rd_block = 0;
    assign fifo_intf_534.fifo_wr_block = 0;
    assign fifo_intf_534.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_534;
    csv_file_dump cstatus_csv_dumper_534;
    df_fifo_monitor fifo_monitor_534;
    df_fifo_intf fifo_intf_535(clock,reset);
    assign fifo_intf_535.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_25_U.if_empty_n;
    assign fifo_intf_535.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_25_U.if_full_n;
    assign fifo_intf_535.fifo_rd_block = 0;
    assign fifo_intf_535.fifo_wr_block = 0;
    assign fifo_intf_535.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_535;
    csv_file_dump cstatus_csv_dumper_535;
    df_fifo_monitor fifo_monitor_535;
    df_fifo_intf fifo_intf_536(clock,reset);
    assign fifo_intf_536.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_25_U.if_empty_n;
    assign fifo_intf_536.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_25_U.if_full_n;
    assign fifo_intf_536.fifo_rd_block = 0;
    assign fifo_intf_536.fifo_wr_block = 0;
    assign fifo_intf_536.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_536;
    csv_file_dump cstatus_csv_dumper_536;
    df_fifo_monitor fifo_monitor_536;
    df_fifo_intf fifo_intf_537(clock,reset);
    assign fifo_intf_537.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_25_U.if_empty_n;
    assign fifo_intf_537.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_25_U.if_full_n;
    assign fifo_intf_537.fifo_rd_block = 0;
    assign fifo_intf_537.fifo_wr_block = 0;
    assign fifo_intf_537.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_537;
    csv_file_dump cstatus_csv_dumper_537;
    df_fifo_monitor fifo_monitor_537;
    df_fifo_intf fifo_intf_538(clock,reset);
    assign fifo_intf_538.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_25_U.if_empty_n;
    assign fifo_intf_538.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_25_U.if_full_n;
    assign fifo_intf_538.fifo_rd_block = 0;
    assign fifo_intf_538.fifo_wr_block = 0;
    assign fifo_intf_538.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_538;
    csv_file_dump cstatus_csv_dumper_538;
    df_fifo_monitor fifo_monitor_538;
    df_fifo_intf fifo_intf_539(clock,reset);
    assign fifo_intf_539.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_25_U.if_empty_n;
    assign fifo_intf_539.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_25_U.if_full_n;
    assign fifo_intf_539.fifo_rd_block = 0;
    assign fifo_intf_539.fifo_wr_block = 0;
    assign fifo_intf_539.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_539;
    csv_file_dump cstatus_csv_dumper_539;
    df_fifo_monitor fifo_monitor_539;
    df_fifo_intf fifo_intf_540(clock,reset);
    assign fifo_intf_540.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_25_U.if_empty_n;
    assign fifo_intf_540.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_25_U.if_full_n;
    assign fifo_intf_540.fifo_rd_block = 0;
    assign fifo_intf_540.fifo_wr_block = 0;
    assign fifo_intf_540.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_540;
    csv_file_dump cstatus_csv_dumper_540;
    df_fifo_monitor fifo_monitor_540;
    df_fifo_intf fifo_intf_541(clock,reset);
    assign fifo_intf_541.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_25_U.if_empty_n;
    assign fifo_intf_541.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_25_U.if_full_n;
    assign fifo_intf_541.fifo_rd_block = 0;
    assign fifo_intf_541.fifo_wr_block = 0;
    assign fifo_intf_541.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_541;
    csv_file_dump cstatus_csv_dumper_541;
    df_fifo_monitor fifo_monitor_541;
    df_fifo_intf fifo_intf_542(clock,reset);
    assign fifo_intf_542.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_25_U.if_empty_n;
    assign fifo_intf_542.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_25_U.if_full_n;
    assign fifo_intf_542.fifo_rd_block = 0;
    assign fifo_intf_542.fifo_wr_block = 0;
    assign fifo_intf_542.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_542;
    csv_file_dump cstatus_csv_dumper_542;
    df_fifo_monitor fifo_monitor_542;
    df_fifo_intf fifo_intf_543(clock,reset);
    assign fifo_intf_543.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_25_U.if_empty_n;
    assign fifo_intf_543.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_25_U.if_full_n;
    assign fifo_intf_543.fifo_rd_block = 0;
    assign fifo_intf_543.fifo_wr_block = 0;
    assign fifo_intf_543.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_543;
    csv_file_dump cstatus_csv_dumper_543;
    df_fifo_monitor fifo_monitor_543;
    df_fifo_intf fifo_intf_544(clock,reset);
    assign fifo_intf_544.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_25_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_25_U.if_empty_n;
    assign fifo_intf_544.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_25_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_25_U.if_full_n;
    assign fifo_intf_544.fifo_rd_block = 0;
    assign fifo_intf_544.fifo_wr_block = 0;
    assign fifo_intf_544.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_544;
    csv_file_dump cstatus_csv_dumper_544;
    df_fifo_monitor fifo_monitor_544;
    df_fifo_intf fifo_intf_545(clock,reset);
    assign fifo_intf_545.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_26_U.if_empty_n;
    assign fifo_intf_545.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_26_U.if_full_n;
    assign fifo_intf_545.fifo_rd_block = 0;
    assign fifo_intf_545.fifo_wr_block = 0;
    assign fifo_intf_545.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_545;
    csv_file_dump cstatus_csv_dumper_545;
    df_fifo_monitor fifo_monitor_545;
    df_fifo_intf fifo_intf_546(clock,reset);
    assign fifo_intf_546.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_26_U.if_empty_n;
    assign fifo_intf_546.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_26_U.if_full_n;
    assign fifo_intf_546.fifo_rd_block = 0;
    assign fifo_intf_546.fifo_wr_block = 0;
    assign fifo_intf_546.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_546;
    csv_file_dump cstatus_csv_dumper_546;
    df_fifo_monitor fifo_monitor_546;
    df_fifo_intf fifo_intf_547(clock,reset);
    assign fifo_intf_547.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_26_U.if_empty_n;
    assign fifo_intf_547.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_26_U.if_full_n;
    assign fifo_intf_547.fifo_rd_block = 0;
    assign fifo_intf_547.fifo_wr_block = 0;
    assign fifo_intf_547.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_547;
    csv_file_dump cstatus_csv_dumper_547;
    df_fifo_monitor fifo_monitor_547;
    df_fifo_intf fifo_intf_548(clock,reset);
    assign fifo_intf_548.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_26_U.if_empty_n;
    assign fifo_intf_548.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_26_U.if_full_n;
    assign fifo_intf_548.fifo_rd_block = 0;
    assign fifo_intf_548.fifo_wr_block = 0;
    assign fifo_intf_548.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_548;
    csv_file_dump cstatus_csv_dumper_548;
    df_fifo_monitor fifo_monitor_548;
    df_fifo_intf fifo_intf_549(clock,reset);
    assign fifo_intf_549.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_26_U.if_empty_n;
    assign fifo_intf_549.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_26_U.if_full_n;
    assign fifo_intf_549.fifo_rd_block = 0;
    assign fifo_intf_549.fifo_wr_block = 0;
    assign fifo_intf_549.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_549;
    csv_file_dump cstatus_csv_dumper_549;
    df_fifo_monitor fifo_monitor_549;
    df_fifo_intf fifo_intf_550(clock,reset);
    assign fifo_intf_550.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_26_U.if_empty_n;
    assign fifo_intf_550.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_26_U.if_full_n;
    assign fifo_intf_550.fifo_rd_block = 0;
    assign fifo_intf_550.fifo_wr_block = 0;
    assign fifo_intf_550.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_550;
    csv_file_dump cstatus_csv_dumper_550;
    df_fifo_monitor fifo_monitor_550;
    df_fifo_intf fifo_intf_551(clock,reset);
    assign fifo_intf_551.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_26_U.if_empty_n;
    assign fifo_intf_551.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_26_U.if_full_n;
    assign fifo_intf_551.fifo_rd_block = 0;
    assign fifo_intf_551.fifo_wr_block = 0;
    assign fifo_intf_551.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_551;
    csv_file_dump cstatus_csv_dumper_551;
    df_fifo_monitor fifo_monitor_551;
    df_fifo_intf fifo_intf_552(clock,reset);
    assign fifo_intf_552.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_26_U.if_empty_n;
    assign fifo_intf_552.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_26_U.if_full_n;
    assign fifo_intf_552.fifo_rd_block = 0;
    assign fifo_intf_552.fifo_wr_block = 0;
    assign fifo_intf_552.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_552;
    csv_file_dump cstatus_csv_dumper_552;
    df_fifo_monitor fifo_monitor_552;
    df_fifo_intf fifo_intf_553(clock,reset);
    assign fifo_intf_553.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_26_U.if_empty_n;
    assign fifo_intf_553.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_26_U.if_full_n;
    assign fifo_intf_553.fifo_rd_block = 0;
    assign fifo_intf_553.fifo_wr_block = 0;
    assign fifo_intf_553.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_553;
    csv_file_dump cstatus_csv_dumper_553;
    df_fifo_monitor fifo_monitor_553;
    df_fifo_intf fifo_intf_554(clock,reset);
    assign fifo_intf_554.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_26_U.if_empty_n;
    assign fifo_intf_554.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_26_U.if_full_n;
    assign fifo_intf_554.fifo_rd_block = 0;
    assign fifo_intf_554.fifo_wr_block = 0;
    assign fifo_intf_554.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_554;
    csv_file_dump cstatus_csv_dumper_554;
    df_fifo_monitor fifo_monitor_554;
    df_fifo_intf fifo_intf_555(clock,reset);
    assign fifo_intf_555.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_26_U.if_empty_n;
    assign fifo_intf_555.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_26_U.if_full_n;
    assign fifo_intf_555.fifo_rd_block = 0;
    assign fifo_intf_555.fifo_wr_block = 0;
    assign fifo_intf_555.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_555;
    csv_file_dump cstatus_csv_dumper_555;
    df_fifo_monitor fifo_monitor_555;
    df_fifo_intf fifo_intf_556(clock,reset);
    assign fifo_intf_556.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_26_U.if_empty_n;
    assign fifo_intf_556.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_26_U.if_full_n;
    assign fifo_intf_556.fifo_rd_block = 0;
    assign fifo_intf_556.fifo_wr_block = 0;
    assign fifo_intf_556.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_556;
    csv_file_dump cstatus_csv_dumper_556;
    df_fifo_monitor fifo_monitor_556;
    df_fifo_intf fifo_intf_557(clock,reset);
    assign fifo_intf_557.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_26_U.if_empty_n;
    assign fifo_intf_557.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_26_U.if_full_n;
    assign fifo_intf_557.fifo_rd_block = 0;
    assign fifo_intf_557.fifo_wr_block = 0;
    assign fifo_intf_557.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_557;
    csv_file_dump cstatus_csv_dumper_557;
    df_fifo_monitor fifo_monitor_557;
    df_fifo_intf fifo_intf_558(clock,reset);
    assign fifo_intf_558.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_26_U.if_empty_n;
    assign fifo_intf_558.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_26_U.if_full_n;
    assign fifo_intf_558.fifo_rd_block = 0;
    assign fifo_intf_558.fifo_wr_block = 0;
    assign fifo_intf_558.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_558;
    csv_file_dump cstatus_csv_dumper_558;
    df_fifo_monitor fifo_monitor_558;
    df_fifo_intf fifo_intf_559(clock,reset);
    assign fifo_intf_559.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_26_U.if_empty_n;
    assign fifo_intf_559.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_26_U.if_full_n;
    assign fifo_intf_559.fifo_rd_block = 0;
    assign fifo_intf_559.fifo_wr_block = 0;
    assign fifo_intf_559.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_559;
    csv_file_dump cstatus_csv_dumper_559;
    df_fifo_monitor fifo_monitor_559;
    df_fifo_intf fifo_intf_560(clock,reset);
    assign fifo_intf_560.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_26_U.if_empty_n;
    assign fifo_intf_560.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_26_U.if_full_n;
    assign fifo_intf_560.fifo_rd_block = 0;
    assign fifo_intf_560.fifo_wr_block = 0;
    assign fifo_intf_560.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_560;
    csv_file_dump cstatus_csv_dumper_560;
    df_fifo_monitor fifo_monitor_560;
    df_fifo_intf fifo_intf_561(clock,reset);
    assign fifo_intf_561.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_26_U.if_empty_n;
    assign fifo_intf_561.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_26_U.if_full_n;
    assign fifo_intf_561.fifo_rd_block = 0;
    assign fifo_intf_561.fifo_wr_block = 0;
    assign fifo_intf_561.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_561;
    csv_file_dump cstatus_csv_dumper_561;
    df_fifo_monitor fifo_monitor_561;
    df_fifo_intf fifo_intf_562(clock,reset);
    assign fifo_intf_562.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_26_U.if_empty_n;
    assign fifo_intf_562.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_26_U.if_full_n;
    assign fifo_intf_562.fifo_rd_block = 0;
    assign fifo_intf_562.fifo_wr_block = 0;
    assign fifo_intf_562.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_562;
    csv_file_dump cstatus_csv_dumper_562;
    df_fifo_monitor fifo_monitor_562;
    df_fifo_intf fifo_intf_563(clock,reset);
    assign fifo_intf_563.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_26_U.if_empty_n;
    assign fifo_intf_563.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_26_U.if_full_n;
    assign fifo_intf_563.fifo_rd_block = 0;
    assign fifo_intf_563.fifo_wr_block = 0;
    assign fifo_intf_563.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_563;
    csv_file_dump cstatus_csv_dumper_563;
    df_fifo_monitor fifo_monitor_563;
    df_fifo_intf fifo_intf_564(clock,reset);
    assign fifo_intf_564.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_26_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_26_U.if_empty_n;
    assign fifo_intf_564.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_26_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_26_U.if_full_n;
    assign fifo_intf_564.fifo_rd_block = 0;
    assign fifo_intf_564.fifo_wr_block = 0;
    assign fifo_intf_564.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_564;
    csv_file_dump cstatus_csv_dumper_564;
    df_fifo_monitor fifo_monitor_564;
    df_fifo_intf fifo_intf_565(clock,reset);
    assign fifo_intf_565.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_27_U.if_empty_n;
    assign fifo_intf_565.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_27_U.if_full_n;
    assign fifo_intf_565.fifo_rd_block = 0;
    assign fifo_intf_565.fifo_wr_block = 0;
    assign fifo_intf_565.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_565;
    csv_file_dump cstatus_csv_dumper_565;
    df_fifo_monitor fifo_monitor_565;
    df_fifo_intf fifo_intf_566(clock,reset);
    assign fifo_intf_566.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_27_U.if_empty_n;
    assign fifo_intf_566.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_27_U.if_full_n;
    assign fifo_intf_566.fifo_rd_block = 0;
    assign fifo_intf_566.fifo_wr_block = 0;
    assign fifo_intf_566.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_566;
    csv_file_dump cstatus_csv_dumper_566;
    df_fifo_monitor fifo_monitor_566;
    df_fifo_intf fifo_intf_567(clock,reset);
    assign fifo_intf_567.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_27_U.if_empty_n;
    assign fifo_intf_567.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_27_U.if_full_n;
    assign fifo_intf_567.fifo_rd_block = 0;
    assign fifo_intf_567.fifo_wr_block = 0;
    assign fifo_intf_567.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_567;
    csv_file_dump cstatus_csv_dumper_567;
    df_fifo_monitor fifo_monitor_567;
    df_fifo_intf fifo_intf_568(clock,reset);
    assign fifo_intf_568.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_27_U.if_empty_n;
    assign fifo_intf_568.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_27_U.if_full_n;
    assign fifo_intf_568.fifo_rd_block = 0;
    assign fifo_intf_568.fifo_wr_block = 0;
    assign fifo_intf_568.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_568;
    csv_file_dump cstatus_csv_dumper_568;
    df_fifo_monitor fifo_monitor_568;
    df_fifo_intf fifo_intf_569(clock,reset);
    assign fifo_intf_569.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_27_U.if_empty_n;
    assign fifo_intf_569.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_27_U.if_full_n;
    assign fifo_intf_569.fifo_rd_block = 0;
    assign fifo_intf_569.fifo_wr_block = 0;
    assign fifo_intf_569.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_569;
    csv_file_dump cstatus_csv_dumper_569;
    df_fifo_monitor fifo_monitor_569;
    df_fifo_intf fifo_intf_570(clock,reset);
    assign fifo_intf_570.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_27_U.if_empty_n;
    assign fifo_intf_570.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_27_U.if_full_n;
    assign fifo_intf_570.fifo_rd_block = 0;
    assign fifo_intf_570.fifo_wr_block = 0;
    assign fifo_intf_570.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_570;
    csv_file_dump cstatus_csv_dumper_570;
    df_fifo_monitor fifo_monitor_570;
    df_fifo_intf fifo_intf_571(clock,reset);
    assign fifo_intf_571.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_27_U.if_empty_n;
    assign fifo_intf_571.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_27_U.if_full_n;
    assign fifo_intf_571.fifo_rd_block = 0;
    assign fifo_intf_571.fifo_wr_block = 0;
    assign fifo_intf_571.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_571;
    csv_file_dump cstatus_csv_dumper_571;
    df_fifo_monitor fifo_monitor_571;
    df_fifo_intf fifo_intf_572(clock,reset);
    assign fifo_intf_572.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_27_U.if_empty_n;
    assign fifo_intf_572.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_27_U.if_full_n;
    assign fifo_intf_572.fifo_rd_block = 0;
    assign fifo_intf_572.fifo_wr_block = 0;
    assign fifo_intf_572.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_572;
    csv_file_dump cstatus_csv_dumper_572;
    df_fifo_monitor fifo_monitor_572;
    df_fifo_intf fifo_intf_573(clock,reset);
    assign fifo_intf_573.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_27_U.if_empty_n;
    assign fifo_intf_573.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_27_U.if_full_n;
    assign fifo_intf_573.fifo_rd_block = 0;
    assign fifo_intf_573.fifo_wr_block = 0;
    assign fifo_intf_573.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_573;
    csv_file_dump cstatus_csv_dumper_573;
    df_fifo_monitor fifo_monitor_573;
    df_fifo_intf fifo_intf_574(clock,reset);
    assign fifo_intf_574.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_27_U.if_empty_n;
    assign fifo_intf_574.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_27_U.if_full_n;
    assign fifo_intf_574.fifo_rd_block = 0;
    assign fifo_intf_574.fifo_wr_block = 0;
    assign fifo_intf_574.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_574;
    csv_file_dump cstatus_csv_dumper_574;
    df_fifo_monitor fifo_monitor_574;
    df_fifo_intf fifo_intf_575(clock,reset);
    assign fifo_intf_575.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_27_U.if_empty_n;
    assign fifo_intf_575.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_27_U.if_full_n;
    assign fifo_intf_575.fifo_rd_block = 0;
    assign fifo_intf_575.fifo_wr_block = 0;
    assign fifo_intf_575.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_575;
    csv_file_dump cstatus_csv_dumper_575;
    df_fifo_monitor fifo_monitor_575;
    df_fifo_intf fifo_intf_576(clock,reset);
    assign fifo_intf_576.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_27_U.if_empty_n;
    assign fifo_intf_576.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_27_U.if_full_n;
    assign fifo_intf_576.fifo_rd_block = 0;
    assign fifo_intf_576.fifo_wr_block = 0;
    assign fifo_intf_576.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_576;
    csv_file_dump cstatus_csv_dumper_576;
    df_fifo_monitor fifo_monitor_576;
    df_fifo_intf fifo_intf_577(clock,reset);
    assign fifo_intf_577.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_27_U.if_empty_n;
    assign fifo_intf_577.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_27_U.if_full_n;
    assign fifo_intf_577.fifo_rd_block = 0;
    assign fifo_intf_577.fifo_wr_block = 0;
    assign fifo_intf_577.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_577;
    csv_file_dump cstatus_csv_dumper_577;
    df_fifo_monitor fifo_monitor_577;
    df_fifo_intf fifo_intf_578(clock,reset);
    assign fifo_intf_578.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_27_U.if_empty_n;
    assign fifo_intf_578.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_27_U.if_full_n;
    assign fifo_intf_578.fifo_rd_block = 0;
    assign fifo_intf_578.fifo_wr_block = 0;
    assign fifo_intf_578.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_578;
    csv_file_dump cstatus_csv_dumper_578;
    df_fifo_monitor fifo_monitor_578;
    df_fifo_intf fifo_intf_579(clock,reset);
    assign fifo_intf_579.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_27_U.if_empty_n;
    assign fifo_intf_579.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_27_U.if_full_n;
    assign fifo_intf_579.fifo_rd_block = 0;
    assign fifo_intf_579.fifo_wr_block = 0;
    assign fifo_intf_579.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_579;
    csv_file_dump cstatus_csv_dumper_579;
    df_fifo_monitor fifo_monitor_579;
    df_fifo_intf fifo_intf_580(clock,reset);
    assign fifo_intf_580.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_27_U.if_empty_n;
    assign fifo_intf_580.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_27_U.if_full_n;
    assign fifo_intf_580.fifo_rd_block = 0;
    assign fifo_intf_580.fifo_wr_block = 0;
    assign fifo_intf_580.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_580;
    csv_file_dump cstatus_csv_dumper_580;
    df_fifo_monitor fifo_monitor_580;
    df_fifo_intf fifo_intf_581(clock,reset);
    assign fifo_intf_581.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_27_U.if_empty_n;
    assign fifo_intf_581.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_27_U.if_full_n;
    assign fifo_intf_581.fifo_rd_block = 0;
    assign fifo_intf_581.fifo_wr_block = 0;
    assign fifo_intf_581.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_581;
    csv_file_dump cstatus_csv_dumper_581;
    df_fifo_monitor fifo_monitor_581;
    df_fifo_intf fifo_intf_582(clock,reset);
    assign fifo_intf_582.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_27_U.if_empty_n;
    assign fifo_intf_582.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_27_U.if_full_n;
    assign fifo_intf_582.fifo_rd_block = 0;
    assign fifo_intf_582.fifo_wr_block = 0;
    assign fifo_intf_582.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_582;
    csv_file_dump cstatus_csv_dumper_582;
    df_fifo_monitor fifo_monitor_582;
    df_fifo_intf fifo_intf_583(clock,reset);
    assign fifo_intf_583.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_27_U.if_empty_n;
    assign fifo_intf_583.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_27_U.if_full_n;
    assign fifo_intf_583.fifo_rd_block = 0;
    assign fifo_intf_583.fifo_wr_block = 0;
    assign fifo_intf_583.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_583;
    csv_file_dump cstatus_csv_dumper_583;
    df_fifo_monitor fifo_monitor_583;
    df_fifo_intf fifo_intf_584(clock,reset);
    assign fifo_intf_584.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_27_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_27_U.if_empty_n;
    assign fifo_intf_584.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_27_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_27_U.if_full_n;
    assign fifo_intf_584.fifo_rd_block = 0;
    assign fifo_intf_584.fifo_wr_block = 0;
    assign fifo_intf_584.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_584;
    csv_file_dump cstatus_csv_dumper_584;
    df_fifo_monitor fifo_monitor_584;
    df_fifo_intf fifo_intf_585(clock,reset);
    assign fifo_intf_585.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_28_U.if_empty_n;
    assign fifo_intf_585.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_28_U.if_full_n;
    assign fifo_intf_585.fifo_rd_block = 0;
    assign fifo_intf_585.fifo_wr_block = 0;
    assign fifo_intf_585.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_585;
    csv_file_dump cstatus_csv_dumper_585;
    df_fifo_monitor fifo_monitor_585;
    df_fifo_intf fifo_intf_586(clock,reset);
    assign fifo_intf_586.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_28_U.if_empty_n;
    assign fifo_intf_586.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_28_U.if_full_n;
    assign fifo_intf_586.fifo_rd_block = 0;
    assign fifo_intf_586.fifo_wr_block = 0;
    assign fifo_intf_586.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_586;
    csv_file_dump cstatus_csv_dumper_586;
    df_fifo_monitor fifo_monitor_586;
    df_fifo_intf fifo_intf_587(clock,reset);
    assign fifo_intf_587.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_28_U.if_empty_n;
    assign fifo_intf_587.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_28_U.if_full_n;
    assign fifo_intf_587.fifo_rd_block = 0;
    assign fifo_intf_587.fifo_wr_block = 0;
    assign fifo_intf_587.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_587;
    csv_file_dump cstatus_csv_dumper_587;
    df_fifo_monitor fifo_monitor_587;
    df_fifo_intf fifo_intf_588(clock,reset);
    assign fifo_intf_588.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_28_U.if_empty_n;
    assign fifo_intf_588.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_28_U.if_full_n;
    assign fifo_intf_588.fifo_rd_block = 0;
    assign fifo_intf_588.fifo_wr_block = 0;
    assign fifo_intf_588.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_588;
    csv_file_dump cstatus_csv_dumper_588;
    df_fifo_monitor fifo_monitor_588;
    df_fifo_intf fifo_intf_589(clock,reset);
    assign fifo_intf_589.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_28_U.if_empty_n;
    assign fifo_intf_589.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_28_U.if_full_n;
    assign fifo_intf_589.fifo_rd_block = 0;
    assign fifo_intf_589.fifo_wr_block = 0;
    assign fifo_intf_589.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_589;
    csv_file_dump cstatus_csv_dumper_589;
    df_fifo_monitor fifo_monitor_589;
    df_fifo_intf fifo_intf_590(clock,reset);
    assign fifo_intf_590.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_28_U.if_empty_n;
    assign fifo_intf_590.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_28_U.if_full_n;
    assign fifo_intf_590.fifo_rd_block = 0;
    assign fifo_intf_590.fifo_wr_block = 0;
    assign fifo_intf_590.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_590;
    csv_file_dump cstatus_csv_dumper_590;
    df_fifo_monitor fifo_monitor_590;
    df_fifo_intf fifo_intf_591(clock,reset);
    assign fifo_intf_591.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_28_U.if_empty_n;
    assign fifo_intf_591.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_28_U.if_full_n;
    assign fifo_intf_591.fifo_rd_block = 0;
    assign fifo_intf_591.fifo_wr_block = 0;
    assign fifo_intf_591.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_591;
    csv_file_dump cstatus_csv_dumper_591;
    df_fifo_monitor fifo_monitor_591;
    df_fifo_intf fifo_intf_592(clock,reset);
    assign fifo_intf_592.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_28_U.if_empty_n;
    assign fifo_intf_592.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_28_U.if_full_n;
    assign fifo_intf_592.fifo_rd_block = 0;
    assign fifo_intf_592.fifo_wr_block = 0;
    assign fifo_intf_592.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_592;
    csv_file_dump cstatus_csv_dumper_592;
    df_fifo_monitor fifo_monitor_592;
    df_fifo_intf fifo_intf_593(clock,reset);
    assign fifo_intf_593.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_28_U.if_empty_n;
    assign fifo_intf_593.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_28_U.if_full_n;
    assign fifo_intf_593.fifo_rd_block = 0;
    assign fifo_intf_593.fifo_wr_block = 0;
    assign fifo_intf_593.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_593;
    csv_file_dump cstatus_csv_dumper_593;
    df_fifo_monitor fifo_monitor_593;
    df_fifo_intf fifo_intf_594(clock,reset);
    assign fifo_intf_594.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_28_U.if_empty_n;
    assign fifo_intf_594.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_28_U.if_full_n;
    assign fifo_intf_594.fifo_rd_block = 0;
    assign fifo_intf_594.fifo_wr_block = 0;
    assign fifo_intf_594.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_594;
    csv_file_dump cstatus_csv_dumper_594;
    df_fifo_monitor fifo_monitor_594;
    df_fifo_intf fifo_intf_595(clock,reset);
    assign fifo_intf_595.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_28_U.if_empty_n;
    assign fifo_intf_595.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_28_U.if_full_n;
    assign fifo_intf_595.fifo_rd_block = 0;
    assign fifo_intf_595.fifo_wr_block = 0;
    assign fifo_intf_595.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_595;
    csv_file_dump cstatus_csv_dumper_595;
    df_fifo_monitor fifo_monitor_595;
    df_fifo_intf fifo_intf_596(clock,reset);
    assign fifo_intf_596.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_28_U.if_empty_n;
    assign fifo_intf_596.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_28_U.if_full_n;
    assign fifo_intf_596.fifo_rd_block = 0;
    assign fifo_intf_596.fifo_wr_block = 0;
    assign fifo_intf_596.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_596;
    csv_file_dump cstatus_csv_dumper_596;
    df_fifo_monitor fifo_monitor_596;
    df_fifo_intf fifo_intf_597(clock,reset);
    assign fifo_intf_597.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_28_U.if_empty_n;
    assign fifo_intf_597.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_28_U.if_full_n;
    assign fifo_intf_597.fifo_rd_block = 0;
    assign fifo_intf_597.fifo_wr_block = 0;
    assign fifo_intf_597.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_597;
    csv_file_dump cstatus_csv_dumper_597;
    df_fifo_monitor fifo_monitor_597;
    df_fifo_intf fifo_intf_598(clock,reset);
    assign fifo_intf_598.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_28_U.if_empty_n;
    assign fifo_intf_598.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_28_U.if_full_n;
    assign fifo_intf_598.fifo_rd_block = 0;
    assign fifo_intf_598.fifo_wr_block = 0;
    assign fifo_intf_598.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_598;
    csv_file_dump cstatus_csv_dumper_598;
    df_fifo_monitor fifo_monitor_598;
    df_fifo_intf fifo_intf_599(clock,reset);
    assign fifo_intf_599.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_28_U.if_empty_n;
    assign fifo_intf_599.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_28_U.if_full_n;
    assign fifo_intf_599.fifo_rd_block = 0;
    assign fifo_intf_599.fifo_wr_block = 0;
    assign fifo_intf_599.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_599;
    csv_file_dump cstatus_csv_dumper_599;
    df_fifo_monitor fifo_monitor_599;
    df_fifo_intf fifo_intf_600(clock,reset);
    assign fifo_intf_600.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_28_U.if_empty_n;
    assign fifo_intf_600.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_28_U.if_full_n;
    assign fifo_intf_600.fifo_rd_block = 0;
    assign fifo_intf_600.fifo_wr_block = 0;
    assign fifo_intf_600.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_600;
    csv_file_dump cstatus_csv_dumper_600;
    df_fifo_monitor fifo_monitor_600;
    df_fifo_intf fifo_intf_601(clock,reset);
    assign fifo_intf_601.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_28_U.if_empty_n;
    assign fifo_intf_601.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_28_U.if_full_n;
    assign fifo_intf_601.fifo_rd_block = 0;
    assign fifo_intf_601.fifo_wr_block = 0;
    assign fifo_intf_601.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_601;
    csv_file_dump cstatus_csv_dumper_601;
    df_fifo_monitor fifo_monitor_601;
    df_fifo_intf fifo_intf_602(clock,reset);
    assign fifo_intf_602.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_28_U.if_empty_n;
    assign fifo_intf_602.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_28_U.if_full_n;
    assign fifo_intf_602.fifo_rd_block = 0;
    assign fifo_intf_602.fifo_wr_block = 0;
    assign fifo_intf_602.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_602;
    csv_file_dump cstatus_csv_dumper_602;
    df_fifo_monitor fifo_monitor_602;
    df_fifo_intf fifo_intf_603(clock,reset);
    assign fifo_intf_603.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_28_U.if_empty_n;
    assign fifo_intf_603.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_28_U.if_full_n;
    assign fifo_intf_603.fifo_rd_block = 0;
    assign fifo_intf_603.fifo_wr_block = 0;
    assign fifo_intf_603.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_603;
    csv_file_dump cstatus_csv_dumper_603;
    df_fifo_monitor fifo_monitor_603;
    df_fifo_intf fifo_intf_604(clock,reset);
    assign fifo_intf_604.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_28_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_28_U.if_empty_n;
    assign fifo_intf_604.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_28_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_28_U.if_full_n;
    assign fifo_intf_604.fifo_rd_block = 0;
    assign fifo_intf_604.fifo_wr_block = 0;
    assign fifo_intf_604.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_604;
    csv_file_dump cstatus_csv_dumper_604;
    df_fifo_monitor fifo_monitor_604;
    df_fifo_intf fifo_intf_605(clock,reset);
    assign fifo_intf_605.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_29_U.if_empty_n;
    assign fifo_intf_605.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_29_U.if_full_n;
    assign fifo_intf_605.fifo_rd_block = 0;
    assign fifo_intf_605.fifo_wr_block = 0;
    assign fifo_intf_605.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_605;
    csv_file_dump cstatus_csv_dumper_605;
    df_fifo_monitor fifo_monitor_605;
    df_fifo_intf fifo_intf_606(clock,reset);
    assign fifo_intf_606.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_29_U.if_empty_n;
    assign fifo_intf_606.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_29_U.if_full_n;
    assign fifo_intf_606.fifo_rd_block = 0;
    assign fifo_intf_606.fifo_wr_block = 0;
    assign fifo_intf_606.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_606;
    csv_file_dump cstatus_csv_dumper_606;
    df_fifo_monitor fifo_monitor_606;
    df_fifo_intf fifo_intf_607(clock,reset);
    assign fifo_intf_607.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_29_U.if_empty_n;
    assign fifo_intf_607.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_29_U.if_full_n;
    assign fifo_intf_607.fifo_rd_block = 0;
    assign fifo_intf_607.fifo_wr_block = 0;
    assign fifo_intf_607.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_607;
    csv_file_dump cstatus_csv_dumper_607;
    df_fifo_monitor fifo_monitor_607;
    df_fifo_intf fifo_intf_608(clock,reset);
    assign fifo_intf_608.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_29_U.if_empty_n;
    assign fifo_intf_608.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_29_U.if_full_n;
    assign fifo_intf_608.fifo_rd_block = 0;
    assign fifo_intf_608.fifo_wr_block = 0;
    assign fifo_intf_608.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_608;
    csv_file_dump cstatus_csv_dumper_608;
    df_fifo_monitor fifo_monitor_608;
    df_fifo_intf fifo_intf_609(clock,reset);
    assign fifo_intf_609.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_29_U.if_empty_n;
    assign fifo_intf_609.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_29_U.if_full_n;
    assign fifo_intf_609.fifo_rd_block = 0;
    assign fifo_intf_609.fifo_wr_block = 0;
    assign fifo_intf_609.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_609;
    csv_file_dump cstatus_csv_dumper_609;
    df_fifo_monitor fifo_monitor_609;
    df_fifo_intf fifo_intf_610(clock,reset);
    assign fifo_intf_610.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_29_U.if_empty_n;
    assign fifo_intf_610.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_29_U.if_full_n;
    assign fifo_intf_610.fifo_rd_block = 0;
    assign fifo_intf_610.fifo_wr_block = 0;
    assign fifo_intf_610.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_610;
    csv_file_dump cstatus_csv_dumper_610;
    df_fifo_monitor fifo_monitor_610;
    df_fifo_intf fifo_intf_611(clock,reset);
    assign fifo_intf_611.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_29_U.if_empty_n;
    assign fifo_intf_611.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_29_U.if_full_n;
    assign fifo_intf_611.fifo_rd_block = 0;
    assign fifo_intf_611.fifo_wr_block = 0;
    assign fifo_intf_611.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_611;
    csv_file_dump cstatus_csv_dumper_611;
    df_fifo_monitor fifo_monitor_611;
    df_fifo_intf fifo_intf_612(clock,reset);
    assign fifo_intf_612.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_29_U.if_empty_n;
    assign fifo_intf_612.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_29_U.if_full_n;
    assign fifo_intf_612.fifo_rd_block = 0;
    assign fifo_intf_612.fifo_wr_block = 0;
    assign fifo_intf_612.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_612;
    csv_file_dump cstatus_csv_dumper_612;
    df_fifo_monitor fifo_monitor_612;
    df_fifo_intf fifo_intf_613(clock,reset);
    assign fifo_intf_613.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_29_U.if_empty_n;
    assign fifo_intf_613.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_29_U.if_full_n;
    assign fifo_intf_613.fifo_rd_block = 0;
    assign fifo_intf_613.fifo_wr_block = 0;
    assign fifo_intf_613.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_613;
    csv_file_dump cstatus_csv_dumper_613;
    df_fifo_monitor fifo_monitor_613;
    df_fifo_intf fifo_intf_614(clock,reset);
    assign fifo_intf_614.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_29_U.if_empty_n;
    assign fifo_intf_614.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_29_U.if_full_n;
    assign fifo_intf_614.fifo_rd_block = 0;
    assign fifo_intf_614.fifo_wr_block = 0;
    assign fifo_intf_614.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_614;
    csv_file_dump cstatus_csv_dumper_614;
    df_fifo_monitor fifo_monitor_614;
    df_fifo_intf fifo_intf_615(clock,reset);
    assign fifo_intf_615.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_29_U.if_empty_n;
    assign fifo_intf_615.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_29_U.if_full_n;
    assign fifo_intf_615.fifo_rd_block = 0;
    assign fifo_intf_615.fifo_wr_block = 0;
    assign fifo_intf_615.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_615;
    csv_file_dump cstatus_csv_dumper_615;
    df_fifo_monitor fifo_monitor_615;
    df_fifo_intf fifo_intf_616(clock,reset);
    assign fifo_intf_616.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_29_U.if_empty_n;
    assign fifo_intf_616.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_29_U.if_full_n;
    assign fifo_intf_616.fifo_rd_block = 0;
    assign fifo_intf_616.fifo_wr_block = 0;
    assign fifo_intf_616.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_616;
    csv_file_dump cstatus_csv_dumper_616;
    df_fifo_monitor fifo_monitor_616;
    df_fifo_intf fifo_intf_617(clock,reset);
    assign fifo_intf_617.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_29_U.if_empty_n;
    assign fifo_intf_617.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_29_U.if_full_n;
    assign fifo_intf_617.fifo_rd_block = 0;
    assign fifo_intf_617.fifo_wr_block = 0;
    assign fifo_intf_617.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_617;
    csv_file_dump cstatus_csv_dumper_617;
    df_fifo_monitor fifo_monitor_617;
    df_fifo_intf fifo_intf_618(clock,reset);
    assign fifo_intf_618.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_29_U.if_empty_n;
    assign fifo_intf_618.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_29_U.if_full_n;
    assign fifo_intf_618.fifo_rd_block = 0;
    assign fifo_intf_618.fifo_wr_block = 0;
    assign fifo_intf_618.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_618;
    csv_file_dump cstatus_csv_dumper_618;
    df_fifo_monitor fifo_monitor_618;
    df_fifo_intf fifo_intf_619(clock,reset);
    assign fifo_intf_619.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_29_U.if_empty_n;
    assign fifo_intf_619.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_29_U.if_full_n;
    assign fifo_intf_619.fifo_rd_block = 0;
    assign fifo_intf_619.fifo_wr_block = 0;
    assign fifo_intf_619.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_619;
    csv_file_dump cstatus_csv_dumper_619;
    df_fifo_monitor fifo_monitor_619;
    df_fifo_intf fifo_intf_620(clock,reset);
    assign fifo_intf_620.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_29_U.if_empty_n;
    assign fifo_intf_620.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_29_U.if_full_n;
    assign fifo_intf_620.fifo_rd_block = 0;
    assign fifo_intf_620.fifo_wr_block = 0;
    assign fifo_intf_620.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_620;
    csv_file_dump cstatus_csv_dumper_620;
    df_fifo_monitor fifo_monitor_620;
    df_fifo_intf fifo_intf_621(clock,reset);
    assign fifo_intf_621.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_29_U.if_empty_n;
    assign fifo_intf_621.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_29_U.if_full_n;
    assign fifo_intf_621.fifo_rd_block = 0;
    assign fifo_intf_621.fifo_wr_block = 0;
    assign fifo_intf_621.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_621;
    csv_file_dump cstatus_csv_dumper_621;
    df_fifo_monitor fifo_monitor_621;
    df_fifo_intf fifo_intf_622(clock,reset);
    assign fifo_intf_622.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_29_U.if_empty_n;
    assign fifo_intf_622.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_29_U.if_full_n;
    assign fifo_intf_622.fifo_rd_block = 0;
    assign fifo_intf_622.fifo_wr_block = 0;
    assign fifo_intf_622.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_622;
    csv_file_dump cstatus_csv_dumper_622;
    df_fifo_monitor fifo_monitor_622;
    df_fifo_intf fifo_intf_623(clock,reset);
    assign fifo_intf_623.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_29_U.if_empty_n;
    assign fifo_intf_623.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_29_U.if_full_n;
    assign fifo_intf_623.fifo_rd_block = 0;
    assign fifo_intf_623.fifo_wr_block = 0;
    assign fifo_intf_623.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_623;
    csv_file_dump cstatus_csv_dumper_623;
    df_fifo_monitor fifo_monitor_623;
    df_fifo_intf fifo_intf_624(clock,reset);
    assign fifo_intf_624.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_29_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_29_U.if_empty_n;
    assign fifo_intf_624.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_29_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_29_U.if_full_n;
    assign fifo_intf_624.fifo_rd_block = 0;
    assign fifo_intf_624.fifo_wr_block = 0;
    assign fifo_intf_624.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_624;
    csv_file_dump cstatus_csv_dumper_624;
    df_fifo_monitor fifo_monitor_624;
    df_fifo_intf fifo_intf_625(clock,reset);
    assign fifo_intf_625.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_30_U.if_empty_n;
    assign fifo_intf_625.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_30_U.if_full_n;
    assign fifo_intf_625.fifo_rd_block = 0;
    assign fifo_intf_625.fifo_wr_block = 0;
    assign fifo_intf_625.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_625;
    csv_file_dump cstatus_csv_dumper_625;
    df_fifo_monitor fifo_monitor_625;
    df_fifo_intf fifo_intf_626(clock,reset);
    assign fifo_intf_626.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_30_U.if_empty_n;
    assign fifo_intf_626.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_30_U.if_full_n;
    assign fifo_intf_626.fifo_rd_block = 0;
    assign fifo_intf_626.fifo_wr_block = 0;
    assign fifo_intf_626.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_626;
    csv_file_dump cstatus_csv_dumper_626;
    df_fifo_monitor fifo_monitor_626;
    df_fifo_intf fifo_intf_627(clock,reset);
    assign fifo_intf_627.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_30_U.if_empty_n;
    assign fifo_intf_627.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_30_U.if_full_n;
    assign fifo_intf_627.fifo_rd_block = 0;
    assign fifo_intf_627.fifo_wr_block = 0;
    assign fifo_intf_627.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_627;
    csv_file_dump cstatus_csv_dumper_627;
    df_fifo_monitor fifo_monitor_627;
    df_fifo_intf fifo_intf_628(clock,reset);
    assign fifo_intf_628.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_30_U.if_empty_n;
    assign fifo_intf_628.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_30_U.if_full_n;
    assign fifo_intf_628.fifo_rd_block = 0;
    assign fifo_intf_628.fifo_wr_block = 0;
    assign fifo_intf_628.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_628;
    csv_file_dump cstatus_csv_dumper_628;
    df_fifo_monitor fifo_monitor_628;
    df_fifo_intf fifo_intf_629(clock,reset);
    assign fifo_intf_629.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_30_U.if_empty_n;
    assign fifo_intf_629.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_30_U.if_full_n;
    assign fifo_intf_629.fifo_rd_block = 0;
    assign fifo_intf_629.fifo_wr_block = 0;
    assign fifo_intf_629.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_629;
    csv_file_dump cstatus_csv_dumper_629;
    df_fifo_monitor fifo_monitor_629;
    df_fifo_intf fifo_intf_630(clock,reset);
    assign fifo_intf_630.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_30_U.if_empty_n;
    assign fifo_intf_630.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_30_U.if_full_n;
    assign fifo_intf_630.fifo_rd_block = 0;
    assign fifo_intf_630.fifo_wr_block = 0;
    assign fifo_intf_630.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_630;
    csv_file_dump cstatus_csv_dumper_630;
    df_fifo_monitor fifo_monitor_630;
    df_fifo_intf fifo_intf_631(clock,reset);
    assign fifo_intf_631.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_30_U.if_empty_n;
    assign fifo_intf_631.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_30_U.if_full_n;
    assign fifo_intf_631.fifo_rd_block = 0;
    assign fifo_intf_631.fifo_wr_block = 0;
    assign fifo_intf_631.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_631;
    csv_file_dump cstatus_csv_dumper_631;
    df_fifo_monitor fifo_monitor_631;
    df_fifo_intf fifo_intf_632(clock,reset);
    assign fifo_intf_632.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_30_U.if_empty_n;
    assign fifo_intf_632.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_30_U.if_full_n;
    assign fifo_intf_632.fifo_rd_block = 0;
    assign fifo_intf_632.fifo_wr_block = 0;
    assign fifo_intf_632.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_632;
    csv_file_dump cstatus_csv_dumper_632;
    df_fifo_monitor fifo_monitor_632;
    df_fifo_intf fifo_intf_633(clock,reset);
    assign fifo_intf_633.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_30_U.if_empty_n;
    assign fifo_intf_633.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_30_U.if_full_n;
    assign fifo_intf_633.fifo_rd_block = 0;
    assign fifo_intf_633.fifo_wr_block = 0;
    assign fifo_intf_633.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_633;
    csv_file_dump cstatus_csv_dumper_633;
    df_fifo_monitor fifo_monitor_633;
    df_fifo_intf fifo_intf_634(clock,reset);
    assign fifo_intf_634.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_30_U.if_empty_n;
    assign fifo_intf_634.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_30_U.if_full_n;
    assign fifo_intf_634.fifo_rd_block = 0;
    assign fifo_intf_634.fifo_wr_block = 0;
    assign fifo_intf_634.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_634;
    csv_file_dump cstatus_csv_dumper_634;
    df_fifo_monitor fifo_monitor_634;
    df_fifo_intf fifo_intf_635(clock,reset);
    assign fifo_intf_635.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_30_U.if_empty_n;
    assign fifo_intf_635.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_30_U.if_full_n;
    assign fifo_intf_635.fifo_rd_block = 0;
    assign fifo_intf_635.fifo_wr_block = 0;
    assign fifo_intf_635.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_635;
    csv_file_dump cstatus_csv_dumper_635;
    df_fifo_monitor fifo_monitor_635;
    df_fifo_intf fifo_intf_636(clock,reset);
    assign fifo_intf_636.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_30_U.if_empty_n;
    assign fifo_intf_636.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_30_U.if_full_n;
    assign fifo_intf_636.fifo_rd_block = 0;
    assign fifo_intf_636.fifo_wr_block = 0;
    assign fifo_intf_636.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_636;
    csv_file_dump cstatus_csv_dumper_636;
    df_fifo_monitor fifo_monitor_636;
    df_fifo_intf fifo_intf_637(clock,reset);
    assign fifo_intf_637.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_30_U.if_empty_n;
    assign fifo_intf_637.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_30_U.if_full_n;
    assign fifo_intf_637.fifo_rd_block = 0;
    assign fifo_intf_637.fifo_wr_block = 0;
    assign fifo_intf_637.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_637;
    csv_file_dump cstatus_csv_dumper_637;
    df_fifo_monitor fifo_monitor_637;
    df_fifo_intf fifo_intf_638(clock,reset);
    assign fifo_intf_638.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_30_U.if_empty_n;
    assign fifo_intf_638.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_30_U.if_full_n;
    assign fifo_intf_638.fifo_rd_block = 0;
    assign fifo_intf_638.fifo_wr_block = 0;
    assign fifo_intf_638.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_638;
    csv_file_dump cstatus_csv_dumper_638;
    df_fifo_monitor fifo_monitor_638;
    df_fifo_intf fifo_intf_639(clock,reset);
    assign fifo_intf_639.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_30_U.if_empty_n;
    assign fifo_intf_639.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_30_U.if_full_n;
    assign fifo_intf_639.fifo_rd_block = 0;
    assign fifo_intf_639.fifo_wr_block = 0;
    assign fifo_intf_639.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_639;
    csv_file_dump cstatus_csv_dumper_639;
    df_fifo_monitor fifo_monitor_639;
    df_fifo_intf fifo_intf_640(clock,reset);
    assign fifo_intf_640.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_30_U.if_empty_n;
    assign fifo_intf_640.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_30_U.if_full_n;
    assign fifo_intf_640.fifo_rd_block = 0;
    assign fifo_intf_640.fifo_wr_block = 0;
    assign fifo_intf_640.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_640;
    csv_file_dump cstatus_csv_dumper_640;
    df_fifo_monitor fifo_monitor_640;
    df_fifo_intf fifo_intf_641(clock,reset);
    assign fifo_intf_641.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_30_U.if_empty_n;
    assign fifo_intf_641.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_30_U.if_full_n;
    assign fifo_intf_641.fifo_rd_block = 0;
    assign fifo_intf_641.fifo_wr_block = 0;
    assign fifo_intf_641.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_641;
    csv_file_dump cstatus_csv_dumper_641;
    df_fifo_monitor fifo_monitor_641;
    df_fifo_intf fifo_intf_642(clock,reset);
    assign fifo_intf_642.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_30_U.if_empty_n;
    assign fifo_intf_642.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_30_U.if_full_n;
    assign fifo_intf_642.fifo_rd_block = 0;
    assign fifo_intf_642.fifo_wr_block = 0;
    assign fifo_intf_642.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_642;
    csv_file_dump cstatus_csv_dumper_642;
    df_fifo_monitor fifo_monitor_642;
    df_fifo_intf fifo_intf_643(clock,reset);
    assign fifo_intf_643.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_30_U.if_empty_n;
    assign fifo_intf_643.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_30_U.if_full_n;
    assign fifo_intf_643.fifo_rd_block = 0;
    assign fifo_intf_643.fifo_wr_block = 0;
    assign fifo_intf_643.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_643;
    csv_file_dump cstatus_csv_dumper_643;
    df_fifo_monitor fifo_monitor_643;
    df_fifo_intf fifo_intf_644(clock,reset);
    assign fifo_intf_644.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_30_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_30_U.if_empty_n;
    assign fifo_intf_644.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_30_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_30_U.if_full_n;
    assign fifo_intf_644.fifo_rd_block = 0;
    assign fifo_intf_644.fifo_wr_block = 0;
    assign fifo_intf_644.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_644;
    csv_file_dump cstatus_csv_dumper_644;
    df_fifo_monitor fifo_monitor_644;
    df_fifo_intf fifo_intf_645(clock,reset);
    assign fifo_intf_645.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_31_U.if_empty_n;
    assign fifo_intf_645.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_31_U.if_full_n;
    assign fifo_intf_645.fifo_rd_block = 0;
    assign fifo_intf_645.fifo_wr_block = 0;
    assign fifo_intf_645.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_645;
    csv_file_dump cstatus_csv_dumper_645;
    df_fifo_monitor fifo_monitor_645;
    df_fifo_intf fifo_intf_646(clock,reset);
    assign fifo_intf_646.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_31_U.if_empty_n;
    assign fifo_intf_646.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_31_U.if_full_n;
    assign fifo_intf_646.fifo_rd_block = 0;
    assign fifo_intf_646.fifo_wr_block = 0;
    assign fifo_intf_646.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_646;
    csv_file_dump cstatus_csv_dumper_646;
    df_fifo_monitor fifo_monitor_646;
    df_fifo_intf fifo_intf_647(clock,reset);
    assign fifo_intf_647.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_31_U.if_empty_n;
    assign fifo_intf_647.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_31_U.if_full_n;
    assign fifo_intf_647.fifo_rd_block = 0;
    assign fifo_intf_647.fifo_wr_block = 0;
    assign fifo_intf_647.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_647;
    csv_file_dump cstatus_csv_dumper_647;
    df_fifo_monitor fifo_monitor_647;
    df_fifo_intf fifo_intf_648(clock,reset);
    assign fifo_intf_648.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_31_U.if_empty_n;
    assign fifo_intf_648.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_31_U.if_full_n;
    assign fifo_intf_648.fifo_rd_block = 0;
    assign fifo_intf_648.fifo_wr_block = 0;
    assign fifo_intf_648.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_648;
    csv_file_dump cstatus_csv_dumper_648;
    df_fifo_monitor fifo_monitor_648;
    df_fifo_intf fifo_intf_649(clock,reset);
    assign fifo_intf_649.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_31_U.if_empty_n;
    assign fifo_intf_649.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_31_U.if_full_n;
    assign fifo_intf_649.fifo_rd_block = 0;
    assign fifo_intf_649.fifo_wr_block = 0;
    assign fifo_intf_649.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_649;
    csv_file_dump cstatus_csv_dumper_649;
    df_fifo_monitor fifo_monitor_649;
    df_fifo_intf fifo_intf_650(clock,reset);
    assign fifo_intf_650.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_31_U.if_empty_n;
    assign fifo_intf_650.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_31_U.if_full_n;
    assign fifo_intf_650.fifo_rd_block = 0;
    assign fifo_intf_650.fifo_wr_block = 0;
    assign fifo_intf_650.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_650;
    csv_file_dump cstatus_csv_dumper_650;
    df_fifo_monitor fifo_monitor_650;
    df_fifo_intf fifo_intf_651(clock,reset);
    assign fifo_intf_651.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_31_U.if_empty_n;
    assign fifo_intf_651.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_31_U.if_full_n;
    assign fifo_intf_651.fifo_rd_block = 0;
    assign fifo_intf_651.fifo_wr_block = 0;
    assign fifo_intf_651.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_651;
    csv_file_dump cstatus_csv_dumper_651;
    df_fifo_monitor fifo_monitor_651;
    df_fifo_intf fifo_intf_652(clock,reset);
    assign fifo_intf_652.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_31_U.if_empty_n;
    assign fifo_intf_652.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_31_U.if_full_n;
    assign fifo_intf_652.fifo_rd_block = 0;
    assign fifo_intf_652.fifo_wr_block = 0;
    assign fifo_intf_652.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_652;
    csv_file_dump cstatus_csv_dumper_652;
    df_fifo_monitor fifo_monitor_652;
    df_fifo_intf fifo_intf_653(clock,reset);
    assign fifo_intf_653.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_31_U.if_empty_n;
    assign fifo_intf_653.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_31_U.if_full_n;
    assign fifo_intf_653.fifo_rd_block = 0;
    assign fifo_intf_653.fifo_wr_block = 0;
    assign fifo_intf_653.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_653;
    csv_file_dump cstatus_csv_dumper_653;
    df_fifo_monitor fifo_monitor_653;
    df_fifo_intf fifo_intf_654(clock,reset);
    assign fifo_intf_654.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_31_U.if_empty_n;
    assign fifo_intf_654.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_31_U.if_full_n;
    assign fifo_intf_654.fifo_rd_block = 0;
    assign fifo_intf_654.fifo_wr_block = 0;
    assign fifo_intf_654.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_654;
    csv_file_dump cstatus_csv_dumper_654;
    df_fifo_monitor fifo_monitor_654;
    df_fifo_intf fifo_intf_655(clock,reset);
    assign fifo_intf_655.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_31_U.if_empty_n;
    assign fifo_intf_655.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_31_U.if_full_n;
    assign fifo_intf_655.fifo_rd_block = 0;
    assign fifo_intf_655.fifo_wr_block = 0;
    assign fifo_intf_655.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_655;
    csv_file_dump cstatus_csv_dumper_655;
    df_fifo_monitor fifo_monitor_655;
    df_fifo_intf fifo_intf_656(clock,reset);
    assign fifo_intf_656.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_31_U.if_empty_n;
    assign fifo_intf_656.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_31_U.if_full_n;
    assign fifo_intf_656.fifo_rd_block = 0;
    assign fifo_intf_656.fifo_wr_block = 0;
    assign fifo_intf_656.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_656;
    csv_file_dump cstatus_csv_dumper_656;
    df_fifo_monitor fifo_monitor_656;
    df_fifo_intf fifo_intf_657(clock,reset);
    assign fifo_intf_657.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_31_U.if_empty_n;
    assign fifo_intf_657.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_31_U.if_full_n;
    assign fifo_intf_657.fifo_rd_block = 0;
    assign fifo_intf_657.fifo_wr_block = 0;
    assign fifo_intf_657.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_657;
    csv_file_dump cstatus_csv_dumper_657;
    df_fifo_monitor fifo_monitor_657;
    df_fifo_intf fifo_intf_658(clock,reset);
    assign fifo_intf_658.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_31_U.if_empty_n;
    assign fifo_intf_658.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_31_U.if_full_n;
    assign fifo_intf_658.fifo_rd_block = 0;
    assign fifo_intf_658.fifo_wr_block = 0;
    assign fifo_intf_658.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_658;
    csv_file_dump cstatus_csv_dumper_658;
    df_fifo_monitor fifo_monitor_658;
    df_fifo_intf fifo_intf_659(clock,reset);
    assign fifo_intf_659.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_31_U.if_empty_n;
    assign fifo_intf_659.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_31_U.if_full_n;
    assign fifo_intf_659.fifo_rd_block = 0;
    assign fifo_intf_659.fifo_wr_block = 0;
    assign fifo_intf_659.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_659;
    csv_file_dump cstatus_csv_dumper_659;
    df_fifo_monitor fifo_monitor_659;
    df_fifo_intf fifo_intf_660(clock,reset);
    assign fifo_intf_660.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_31_U.if_empty_n;
    assign fifo_intf_660.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_31_U.if_full_n;
    assign fifo_intf_660.fifo_rd_block = 0;
    assign fifo_intf_660.fifo_wr_block = 0;
    assign fifo_intf_660.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_660;
    csv_file_dump cstatus_csv_dumper_660;
    df_fifo_monitor fifo_monitor_660;
    df_fifo_intf fifo_intf_661(clock,reset);
    assign fifo_intf_661.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_31_U.if_empty_n;
    assign fifo_intf_661.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_31_U.if_full_n;
    assign fifo_intf_661.fifo_rd_block = 0;
    assign fifo_intf_661.fifo_wr_block = 0;
    assign fifo_intf_661.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_661;
    csv_file_dump cstatus_csv_dumper_661;
    df_fifo_monitor fifo_monitor_661;
    df_fifo_intf fifo_intf_662(clock,reset);
    assign fifo_intf_662.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_31_U.if_empty_n;
    assign fifo_intf_662.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_31_U.if_full_n;
    assign fifo_intf_662.fifo_rd_block = 0;
    assign fifo_intf_662.fifo_wr_block = 0;
    assign fifo_intf_662.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_662;
    csv_file_dump cstatus_csv_dumper_662;
    df_fifo_monitor fifo_monitor_662;
    df_fifo_intf fifo_intf_663(clock,reset);
    assign fifo_intf_663.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_31_U.if_empty_n;
    assign fifo_intf_663.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_31_U.if_full_n;
    assign fifo_intf_663.fifo_rd_block = 0;
    assign fifo_intf_663.fifo_wr_block = 0;
    assign fifo_intf_663.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_663;
    csv_file_dump cstatus_csv_dumper_663;
    df_fifo_monitor fifo_monitor_663;
    df_fifo_intf fifo_intf_664(clock,reset);
    assign fifo_intf_664.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_31_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_31_U.if_empty_n;
    assign fifo_intf_664.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_31_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_31_U.if_full_n;
    assign fifo_intf_664.fifo_rd_block = 0;
    assign fifo_intf_664.fifo_wr_block = 0;
    assign fifo_intf_664.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_664;
    csv_file_dump cstatus_csv_dumper_664;
    df_fifo_monitor fifo_monitor_664;
    df_fifo_intf fifo_intf_665(clock,reset);
    assign fifo_intf_665.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_32_U.if_empty_n;
    assign fifo_intf_665.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_32_U.if_full_n;
    assign fifo_intf_665.fifo_rd_block = 0;
    assign fifo_intf_665.fifo_wr_block = 0;
    assign fifo_intf_665.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_665;
    csv_file_dump cstatus_csv_dumper_665;
    df_fifo_monitor fifo_monitor_665;
    df_fifo_intf fifo_intf_666(clock,reset);
    assign fifo_intf_666.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_32_U.if_empty_n;
    assign fifo_intf_666.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_32_U.if_full_n;
    assign fifo_intf_666.fifo_rd_block = 0;
    assign fifo_intf_666.fifo_wr_block = 0;
    assign fifo_intf_666.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_666;
    csv_file_dump cstatus_csv_dumper_666;
    df_fifo_monitor fifo_monitor_666;
    df_fifo_intf fifo_intf_667(clock,reset);
    assign fifo_intf_667.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_32_U.if_empty_n;
    assign fifo_intf_667.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_32_U.if_full_n;
    assign fifo_intf_667.fifo_rd_block = 0;
    assign fifo_intf_667.fifo_wr_block = 0;
    assign fifo_intf_667.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_667;
    csv_file_dump cstatus_csv_dumper_667;
    df_fifo_monitor fifo_monitor_667;
    df_fifo_intf fifo_intf_668(clock,reset);
    assign fifo_intf_668.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_32_U.if_empty_n;
    assign fifo_intf_668.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_32_U.if_full_n;
    assign fifo_intf_668.fifo_rd_block = 0;
    assign fifo_intf_668.fifo_wr_block = 0;
    assign fifo_intf_668.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_668;
    csv_file_dump cstatus_csv_dumper_668;
    df_fifo_monitor fifo_monitor_668;
    df_fifo_intf fifo_intf_669(clock,reset);
    assign fifo_intf_669.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_32_U.if_empty_n;
    assign fifo_intf_669.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_32_U.if_full_n;
    assign fifo_intf_669.fifo_rd_block = 0;
    assign fifo_intf_669.fifo_wr_block = 0;
    assign fifo_intf_669.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_669;
    csv_file_dump cstatus_csv_dumper_669;
    df_fifo_monitor fifo_monitor_669;
    df_fifo_intf fifo_intf_670(clock,reset);
    assign fifo_intf_670.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_32_U.if_empty_n;
    assign fifo_intf_670.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_32_U.if_full_n;
    assign fifo_intf_670.fifo_rd_block = 0;
    assign fifo_intf_670.fifo_wr_block = 0;
    assign fifo_intf_670.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_670;
    csv_file_dump cstatus_csv_dumper_670;
    df_fifo_monitor fifo_monitor_670;
    df_fifo_intf fifo_intf_671(clock,reset);
    assign fifo_intf_671.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_32_U.if_empty_n;
    assign fifo_intf_671.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_32_U.if_full_n;
    assign fifo_intf_671.fifo_rd_block = 0;
    assign fifo_intf_671.fifo_wr_block = 0;
    assign fifo_intf_671.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_671;
    csv_file_dump cstatus_csv_dumper_671;
    df_fifo_monitor fifo_monitor_671;
    df_fifo_intf fifo_intf_672(clock,reset);
    assign fifo_intf_672.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_32_U.if_empty_n;
    assign fifo_intf_672.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_32_U.if_full_n;
    assign fifo_intf_672.fifo_rd_block = 0;
    assign fifo_intf_672.fifo_wr_block = 0;
    assign fifo_intf_672.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_672;
    csv_file_dump cstatus_csv_dumper_672;
    df_fifo_monitor fifo_monitor_672;
    df_fifo_intf fifo_intf_673(clock,reset);
    assign fifo_intf_673.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_32_U.if_empty_n;
    assign fifo_intf_673.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_32_U.if_full_n;
    assign fifo_intf_673.fifo_rd_block = 0;
    assign fifo_intf_673.fifo_wr_block = 0;
    assign fifo_intf_673.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_673;
    csv_file_dump cstatus_csv_dumper_673;
    df_fifo_monitor fifo_monitor_673;
    df_fifo_intf fifo_intf_674(clock,reset);
    assign fifo_intf_674.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_32_U.if_empty_n;
    assign fifo_intf_674.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_32_U.if_full_n;
    assign fifo_intf_674.fifo_rd_block = 0;
    assign fifo_intf_674.fifo_wr_block = 0;
    assign fifo_intf_674.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_674;
    csv_file_dump cstatus_csv_dumper_674;
    df_fifo_monitor fifo_monitor_674;
    df_fifo_intf fifo_intf_675(clock,reset);
    assign fifo_intf_675.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_32_U.if_empty_n;
    assign fifo_intf_675.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_32_U.if_full_n;
    assign fifo_intf_675.fifo_rd_block = 0;
    assign fifo_intf_675.fifo_wr_block = 0;
    assign fifo_intf_675.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_675;
    csv_file_dump cstatus_csv_dumper_675;
    df_fifo_monitor fifo_monitor_675;
    df_fifo_intf fifo_intf_676(clock,reset);
    assign fifo_intf_676.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_32_U.if_empty_n;
    assign fifo_intf_676.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_32_U.if_full_n;
    assign fifo_intf_676.fifo_rd_block = 0;
    assign fifo_intf_676.fifo_wr_block = 0;
    assign fifo_intf_676.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_676;
    csv_file_dump cstatus_csv_dumper_676;
    df_fifo_monitor fifo_monitor_676;
    df_fifo_intf fifo_intf_677(clock,reset);
    assign fifo_intf_677.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_32_U.if_empty_n;
    assign fifo_intf_677.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_32_U.if_full_n;
    assign fifo_intf_677.fifo_rd_block = 0;
    assign fifo_intf_677.fifo_wr_block = 0;
    assign fifo_intf_677.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_677;
    csv_file_dump cstatus_csv_dumper_677;
    df_fifo_monitor fifo_monitor_677;
    df_fifo_intf fifo_intf_678(clock,reset);
    assign fifo_intf_678.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_32_U.if_empty_n;
    assign fifo_intf_678.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_32_U.if_full_n;
    assign fifo_intf_678.fifo_rd_block = 0;
    assign fifo_intf_678.fifo_wr_block = 0;
    assign fifo_intf_678.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_678;
    csv_file_dump cstatus_csv_dumper_678;
    df_fifo_monitor fifo_monitor_678;
    df_fifo_intf fifo_intf_679(clock,reset);
    assign fifo_intf_679.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_32_U.if_empty_n;
    assign fifo_intf_679.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_32_U.if_full_n;
    assign fifo_intf_679.fifo_rd_block = 0;
    assign fifo_intf_679.fifo_wr_block = 0;
    assign fifo_intf_679.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_679;
    csv_file_dump cstatus_csv_dumper_679;
    df_fifo_monitor fifo_monitor_679;
    df_fifo_intf fifo_intf_680(clock,reset);
    assign fifo_intf_680.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_32_U.if_empty_n;
    assign fifo_intf_680.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_32_U.if_full_n;
    assign fifo_intf_680.fifo_rd_block = 0;
    assign fifo_intf_680.fifo_wr_block = 0;
    assign fifo_intf_680.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_680;
    csv_file_dump cstatus_csv_dumper_680;
    df_fifo_monitor fifo_monitor_680;
    df_fifo_intf fifo_intf_681(clock,reset);
    assign fifo_intf_681.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_32_U.if_empty_n;
    assign fifo_intf_681.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_32_U.if_full_n;
    assign fifo_intf_681.fifo_rd_block = 0;
    assign fifo_intf_681.fifo_wr_block = 0;
    assign fifo_intf_681.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_681;
    csv_file_dump cstatus_csv_dumper_681;
    df_fifo_monitor fifo_monitor_681;
    df_fifo_intf fifo_intf_682(clock,reset);
    assign fifo_intf_682.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_32_U.if_empty_n;
    assign fifo_intf_682.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_32_U.if_full_n;
    assign fifo_intf_682.fifo_rd_block = 0;
    assign fifo_intf_682.fifo_wr_block = 0;
    assign fifo_intf_682.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_682;
    csv_file_dump cstatus_csv_dumper_682;
    df_fifo_monitor fifo_monitor_682;
    df_fifo_intf fifo_intf_683(clock,reset);
    assign fifo_intf_683.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_32_U.if_empty_n;
    assign fifo_intf_683.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_32_U.if_full_n;
    assign fifo_intf_683.fifo_rd_block = 0;
    assign fifo_intf_683.fifo_wr_block = 0;
    assign fifo_intf_683.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_683;
    csv_file_dump cstatus_csv_dumper_683;
    df_fifo_monitor fifo_monitor_683;
    df_fifo_intf fifo_intf_684(clock,reset);
    assign fifo_intf_684.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_32_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_32_U.if_empty_n;
    assign fifo_intf_684.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_32_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_32_U.if_full_n;
    assign fifo_intf_684.fifo_rd_block = 0;
    assign fifo_intf_684.fifo_wr_block = 0;
    assign fifo_intf_684.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_684;
    csv_file_dump cstatus_csv_dumper_684;
    df_fifo_monitor fifo_monitor_684;
    df_fifo_intf fifo_intf_685(clock,reset);
    assign fifo_intf_685.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_33_U.if_empty_n;
    assign fifo_intf_685.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_33_U.if_full_n;
    assign fifo_intf_685.fifo_rd_block = 0;
    assign fifo_intf_685.fifo_wr_block = 0;
    assign fifo_intf_685.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_685;
    csv_file_dump cstatus_csv_dumper_685;
    df_fifo_monitor fifo_monitor_685;
    df_fifo_intf fifo_intf_686(clock,reset);
    assign fifo_intf_686.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_33_U.if_empty_n;
    assign fifo_intf_686.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_33_U.if_full_n;
    assign fifo_intf_686.fifo_rd_block = 0;
    assign fifo_intf_686.fifo_wr_block = 0;
    assign fifo_intf_686.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_686;
    csv_file_dump cstatus_csv_dumper_686;
    df_fifo_monitor fifo_monitor_686;
    df_fifo_intf fifo_intf_687(clock,reset);
    assign fifo_intf_687.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_33_U.if_empty_n;
    assign fifo_intf_687.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_33_U.if_full_n;
    assign fifo_intf_687.fifo_rd_block = 0;
    assign fifo_intf_687.fifo_wr_block = 0;
    assign fifo_intf_687.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_687;
    csv_file_dump cstatus_csv_dumper_687;
    df_fifo_monitor fifo_monitor_687;
    df_fifo_intf fifo_intf_688(clock,reset);
    assign fifo_intf_688.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_33_U.if_empty_n;
    assign fifo_intf_688.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_33_U.if_full_n;
    assign fifo_intf_688.fifo_rd_block = 0;
    assign fifo_intf_688.fifo_wr_block = 0;
    assign fifo_intf_688.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_688;
    csv_file_dump cstatus_csv_dumper_688;
    df_fifo_monitor fifo_monitor_688;
    df_fifo_intf fifo_intf_689(clock,reset);
    assign fifo_intf_689.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_33_U.if_empty_n;
    assign fifo_intf_689.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_33_U.if_full_n;
    assign fifo_intf_689.fifo_rd_block = 0;
    assign fifo_intf_689.fifo_wr_block = 0;
    assign fifo_intf_689.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_689;
    csv_file_dump cstatus_csv_dumper_689;
    df_fifo_monitor fifo_monitor_689;
    df_fifo_intf fifo_intf_690(clock,reset);
    assign fifo_intf_690.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_33_U.if_empty_n;
    assign fifo_intf_690.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_33_U.if_full_n;
    assign fifo_intf_690.fifo_rd_block = 0;
    assign fifo_intf_690.fifo_wr_block = 0;
    assign fifo_intf_690.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_690;
    csv_file_dump cstatus_csv_dumper_690;
    df_fifo_monitor fifo_monitor_690;
    df_fifo_intf fifo_intf_691(clock,reset);
    assign fifo_intf_691.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_33_U.if_empty_n;
    assign fifo_intf_691.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_33_U.if_full_n;
    assign fifo_intf_691.fifo_rd_block = 0;
    assign fifo_intf_691.fifo_wr_block = 0;
    assign fifo_intf_691.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_691;
    csv_file_dump cstatus_csv_dumper_691;
    df_fifo_monitor fifo_monitor_691;
    df_fifo_intf fifo_intf_692(clock,reset);
    assign fifo_intf_692.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_33_U.if_empty_n;
    assign fifo_intf_692.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_33_U.if_full_n;
    assign fifo_intf_692.fifo_rd_block = 0;
    assign fifo_intf_692.fifo_wr_block = 0;
    assign fifo_intf_692.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_692;
    csv_file_dump cstatus_csv_dumper_692;
    df_fifo_monitor fifo_monitor_692;
    df_fifo_intf fifo_intf_693(clock,reset);
    assign fifo_intf_693.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_33_U.if_empty_n;
    assign fifo_intf_693.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_33_U.if_full_n;
    assign fifo_intf_693.fifo_rd_block = 0;
    assign fifo_intf_693.fifo_wr_block = 0;
    assign fifo_intf_693.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_693;
    csv_file_dump cstatus_csv_dumper_693;
    df_fifo_monitor fifo_monitor_693;
    df_fifo_intf fifo_intf_694(clock,reset);
    assign fifo_intf_694.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_33_U.if_empty_n;
    assign fifo_intf_694.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_33_U.if_full_n;
    assign fifo_intf_694.fifo_rd_block = 0;
    assign fifo_intf_694.fifo_wr_block = 0;
    assign fifo_intf_694.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_694;
    csv_file_dump cstatus_csv_dumper_694;
    df_fifo_monitor fifo_monitor_694;
    df_fifo_intf fifo_intf_695(clock,reset);
    assign fifo_intf_695.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_33_U.if_empty_n;
    assign fifo_intf_695.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_33_U.if_full_n;
    assign fifo_intf_695.fifo_rd_block = 0;
    assign fifo_intf_695.fifo_wr_block = 0;
    assign fifo_intf_695.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_695;
    csv_file_dump cstatus_csv_dumper_695;
    df_fifo_monitor fifo_monitor_695;
    df_fifo_intf fifo_intf_696(clock,reset);
    assign fifo_intf_696.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_33_U.if_empty_n;
    assign fifo_intf_696.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_33_U.if_full_n;
    assign fifo_intf_696.fifo_rd_block = 0;
    assign fifo_intf_696.fifo_wr_block = 0;
    assign fifo_intf_696.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_696;
    csv_file_dump cstatus_csv_dumper_696;
    df_fifo_monitor fifo_monitor_696;
    df_fifo_intf fifo_intf_697(clock,reset);
    assign fifo_intf_697.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_33_U.if_empty_n;
    assign fifo_intf_697.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_33_U.if_full_n;
    assign fifo_intf_697.fifo_rd_block = 0;
    assign fifo_intf_697.fifo_wr_block = 0;
    assign fifo_intf_697.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_697;
    csv_file_dump cstatus_csv_dumper_697;
    df_fifo_monitor fifo_monitor_697;
    df_fifo_intf fifo_intf_698(clock,reset);
    assign fifo_intf_698.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_33_U.if_empty_n;
    assign fifo_intf_698.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_33_U.if_full_n;
    assign fifo_intf_698.fifo_rd_block = 0;
    assign fifo_intf_698.fifo_wr_block = 0;
    assign fifo_intf_698.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_698;
    csv_file_dump cstatus_csv_dumper_698;
    df_fifo_monitor fifo_monitor_698;
    df_fifo_intf fifo_intf_699(clock,reset);
    assign fifo_intf_699.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_33_U.if_empty_n;
    assign fifo_intf_699.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_33_U.if_full_n;
    assign fifo_intf_699.fifo_rd_block = 0;
    assign fifo_intf_699.fifo_wr_block = 0;
    assign fifo_intf_699.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_699;
    csv_file_dump cstatus_csv_dumper_699;
    df_fifo_monitor fifo_monitor_699;
    df_fifo_intf fifo_intf_700(clock,reset);
    assign fifo_intf_700.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_33_U.if_empty_n;
    assign fifo_intf_700.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_33_U.if_full_n;
    assign fifo_intf_700.fifo_rd_block = 0;
    assign fifo_intf_700.fifo_wr_block = 0;
    assign fifo_intf_700.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_700;
    csv_file_dump cstatus_csv_dumper_700;
    df_fifo_monitor fifo_monitor_700;
    df_fifo_intf fifo_intf_701(clock,reset);
    assign fifo_intf_701.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_33_U.if_empty_n;
    assign fifo_intf_701.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_33_U.if_full_n;
    assign fifo_intf_701.fifo_rd_block = 0;
    assign fifo_intf_701.fifo_wr_block = 0;
    assign fifo_intf_701.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_701;
    csv_file_dump cstatus_csv_dumper_701;
    df_fifo_monitor fifo_monitor_701;
    df_fifo_intf fifo_intf_702(clock,reset);
    assign fifo_intf_702.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_33_U.if_empty_n;
    assign fifo_intf_702.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_33_U.if_full_n;
    assign fifo_intf_702.fifo_rd_block = 0;
    assign fifo_intf_702.fifo_wr_block = 0;
    assign fifo_intf_702.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_702;
    csv_file_dump cstatus_csv_dumper_702;
    df_fifo_monitor fifo_monitor_702;
    df_fifo_intf fifo_intf_703(clock,reset);
    assign fifo_intf_703.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_33_U.if_empty_n;
    assign fifo_intf_703.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_33_U.if_full_n;
    assign fifo_intf_703.fifo_rd_block = 0;
    assign fifo_intf_703.fifo_wr_block = 0;
    assign fifo_intf_703.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_703;
    csv_file_dump cstatus_csv_dumper_703;
    df_fifo_monitor fifo_monitor_703;
    df_fifo_intf fifo_intf_704(clock,reset);
    assign fifo_intf_704.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_33_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_33_U.if_empty_n;
    assign fifo_intf_704.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_33_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_33_U.if_full_n;
    assign fifo_intf_704.fifo_rd_block = 0;
    assign fifo_intf_704.fifo_wr_block = 0;
    assign fifo_intf_704.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_704;
    csv_file_dump cstatus_csv_dumper_704;
    df_fifo_monitor fifo_monitor_704;
    df_fifo_intf fifo_intf_705(clock,reset);
    assign fifo_intf_705.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_34_U.if_empty_n;
    assign fifo_intf_705.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_34_U.if_full_n;
    assign fifo_intf_705.fifo_rd_block = 0;
    assign fifo_intf_705.fifo_wr_block = 0;
    assign fifo_intf_705.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_705;
    csv_file_dump cstatus_csv_dumper_705;
    df_fifo_monitor fifo_monitor_705;
    df_fifo_intf fifo_intf_706(clock,reset);
    assign fifo_intf_706.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_34_U.if_empty_n;
    assign fifo_intf_706.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_34_U.if_full_n;
    assign fifo_intf_706.fifo_rd_block = 0;
    assign fifo_intf_706.fifo_wr_block = 0;
    assign fifo_intf_706.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_706;
    csv_file_dump cstatus_csv_dumper_706;
    df_fifo_monitor fifo_monitor_706;
    df_fifo_intf fifo_intf_707(clock,reset);
    assign fifo_intf_707.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_34_U.if_empty_n;
    assign fifo_intf_707.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_34_U.if_full_n;
    assign fifo_intf_707.fifo_rd_block = 0;
    assign fifo_intf_707.fifo_wr_block = 0;
    assign fifo_intf_707.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_707;
    csv_file_dump cstatus_csv_dumper_707;
    df_fifo_monitor fifo_monitor_707;
    df_fifo_intf fifo_intf_708(clock,reset);
    assign fifo_intf_708.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_34_U.if_empty_n;
    assign fifo_intf_708.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_34_U.if_full_n;
    assign fifo_intf_708.fifo_rd_block = 0;
    assign fifo_intf_708.fifo_wr_block = 0;
    assign fifo_intf_708.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_708;
    csv_file_dump cstatus_csv_dumper_708;
    df_fifo_monitor fifo_monitor_708;
    df_fifo_intf fifo_intf_709(clock,reset);
    assign fifo_intf_709.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_34_U.if_empty_n;
    assign fifo_intf_709.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_34_U.if_full_n;
    assign fifo_intf_709.fifo_rd_block = 0;
    assign fifo_intf_709.fifo_wr_block = 0;
    assign fifo_intf_709.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_709;
    csv_file_dump cstatus_csv_dumper_709;
    df_fifo_monitor fifo_monitor_709;
    df_fifo_intf fifo_intf_710(clock,reset);
    assign fifo_intf_710.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_34_U.if_empty_n;
    assign fifo_intf_710.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_34_U.if_full_n;
    assign fifo_intf_710.fifo_rd_block = 0;
    assign fifo_intf_710.fifo_wr_block = 0;
    assign fifo_intf_710.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_710;
    csv_file_dump cstatus_csv_dumper_710;
    df_fifo_monitor fifo_monitor_710;
    df_fifo_intf fifo_intf_711(clock,reset);
    assign fifo_intf_711.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_34_U.if_empty_n;
    assign fifo_intf_711.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_34_U.if_full_n;
    assign fifo_intf_711.fifo_rd_block = 0;
    assign fifo_intf_711.fifo_wr_block = 0;
    assign fifo_intf_711.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_711;
    csv_file_dump cstatus_csv_dumper_711;
    df_fifo_monitor fifo_monitor_711;
    df_fifo_intf fifo_intf_712(clock,reset);
    assign fifo_intf_712.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_34_U.if_empty_n;
    assign fifo_intf_712.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_34_U.if_full_n;
    assign fifo_intf_712.fifo_rd_block = 0;
    assign fifo_intf_712.fifo_wr_block = 0;
    assign fifo_intf_712.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_712;
    csv_file_dump cstatus_csv_dumper_712;
    df_fifo_monitor fifo_monitor_712;
    df_fifo_intf fifo_intf_713(clock,reset);
    assign fifo_intf_713.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_34_U.if_empty_n;
    assign fifo_intf_713.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_34_U.if_full_n;
    assign fifo_intf_713.fifo_rd_block = 0;
    assign fifo_intf_713.fifo_wr_block = 0;
    assign fifo_intf_713.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_713;
    csv_file_dump cstatus_csv_dumper_713;
    df_fifo_monitor fifo_monitor_713;
    df_fifo_intf fifo_intf_714(clock,reset);
    assign fifo_intf_714.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_34_U.if_empty_n;
    assign fifo_intf_714.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_34_U.if_full_n;
    assign fifo_intf_714.fifo_rd_block = 0;
    assign fifo_intf_714.fifo_wr_block = 0;
    assign fifo_intf_714.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_714;
    csv_file_dump cstatus_csv_dumper_714;
    df_fifo_monitor fifo_monitor_714;
    df_fifo_intf fifo_intf_715(clock,reset);
    assign fifo_intf_715.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_34_U.if_empty_n;
    assign fifo_intf_715.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_34_U.if_full_n;
    assign fifo_intf_715.fifo_rd_block = 0;
    assign fifo_intf_715.fifo_wr_block = 0;
    assign fifo_intf_715.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_715;
    csv_file_dump cstatus_csv_dumper_715;
    df_fifo_monitor fifo_monitor_715;
    df_fifo_intf fifo_intf_716(clock,reset);
    assign fifo_intf_716.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_34_U.if_empty_n;
    assign fifo_intf_716.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_34_U.if_full_n;
    assign fifo_intf_716.fifo_rd_block = 0;
    assign fifo_intf_716.fifo_wr_block = 0;
    assign fifo_intf_716.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_716;
    csv_file_dump cstatus_csv_dumper_716;
    df_fifo_monitor fifo_monitor_716;
    df_fifo_intf fifo_intf_717(clock,reset);
    assign fifo_intf_717.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_34_U.if_empty_n;
    assign fifo_intf_717.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_34_U.if_full_n;
    assign fifo_intf_717.fifo_rd_block = 0;
    assign fifo_intf_717.fifo_wr_block = 0;
    assign fifo_intf_717.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_717;
    csv_file_dump cstatus_csv_dumper_717;
    df_fifo_monitor fifo_monitor_717;
    df_fifo_intf fifo_intf_718(clock,reset);
    assign fifo_intf_718.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_34_U.if_empty_n;
    assign fifo_intf_718.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_34_U.if_full_n;
    assign fifo_intf_718.fifo_rd_block = 0;
    assign fifo_intf_718.fifo_wr_block = 0;
    assign fifo_intf_718.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_718;
    csv_file_dump cstatus_csv_dumper_718;
    df_fifo_monitor fifo_monitor_718;
    df_fifo_intf fifo_intf_719(clock,reset);
    assign fifo_intf_719.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_34_U.if_empty_n;
    assign fifo_intf_719.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_34_U.if_full_n;
    assign fifo_intf_719.fifo_rd_block = 0;
    assign fifo_intf_719.fifo_wr_block = 0;
    assign fifo_intf_719.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_719;
    csv_file_dump cstatus_csv_dumper_719;
    df_fifo_monitor fifo_monitor_719;
    df_fifo_intf fifo_intf_720(clock,reset);
    assign fifo_intf_720.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_34_U.if_empty_n;
    assign fifo_intf_720.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_34_U.if_full_n;
    assign fifo_intf_720.fifo_rd_block = 0;
    assign fifo_intf_720.fifo_wr_block = 0;
    assign fifo_intf_720.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_720;
    csv_file_dump cstatus_csv_dumper_720;
    df_fifo_monitor fifo_monitor_720;
    df_fifo_intf fifo_intf_721(clock,reset);
    assign fifo_intf_721.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_34_U.if_empty_n;
    assign fifo_intf_721.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_34_U.if_full_n;
    assign fifo_intf_721.fifo_rd_block = 0;
    assign fifo_intf_721.fifo_wr_block = 0;
    assign fifo_intf_721.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_721;
    csv_file_dump cstatus_csv_dumper_721;
    df_fifo_monitor fifo_monitor_721;
    df_fifo_intf fifo_intf_722(clock,reset);
    assign fifo_intf_722.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_34_U.if_empty_n;
    assign fifo_intf_722.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_34_U.if_full_n;
    assign fifo_intf_722.fifo_rd_block = 0;
    assign fifo_intf_722.fifo_wr_block = 0;
    assign fifo_intf_722.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_722;
    csv_file_dump cstatus_csv_dumper_722;
    df_fifo_monitor fifo_monitor_722;
    df_fifo_intf fifo_intf_723(clock,reset);
    assign fifo_intf_723.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_34_U.if_empty_n;
    assign fifo_intf_723.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_34_U.if_full_n;
    assign fifo_intf_723.fifo_rd_block = 0;
    assign fifo_intf_723.fifo_wr_block = 0;
    assign fifo_intf_723.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_723;
    csv_file_dump cstatus_csv_dumper_723;
    df_fifo_monitor fifo_monitor_723;
    df_fifo_intf fifo_intf_724(clock,reset);
    assign fifo_intf_724.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_34_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_34_U.if_empty_n;
    assign fifo_intf_724.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_34_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_34_U.if_full_n;
    assign fifo_intf_724.fifo_rd_block = 0;
    assign fifo_intf_724.fifo_wr_block = 0;
    assign fifo_intf_724.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_724;
    csv_file_dump cstatus_csv_dumper_724;
    df_fifo_monitor fifo_monitor_724;
    df_fifo_intf fifo_intf_725(clock,reset);
    assign fifo_intf_725.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_35_U.if_empty_n;
    assign fifo_intf_725.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_35_U.if_full_n;
    assign fifo_intf_725.fifo_rd_block = 0;
    assign fifo_intf_725.fifo_wr_block = 0;
    assign fifo_intf_725.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_725;
    csv_file_dump cstatus_csv_dumper_725;
    df_fifo_monitor fifo_monitor_725;
    df_fifo_intf fifo_intf_726(clock,reset);
    assign fifo_intf_726.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_35_U.if_empty_n;
    assign fifo_intf_726.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_35_U.if_full_n;
    assign fifo_intf_726.fifo_rd_block = 0;
    assign fifo_intf_726.fifo_wr_block = 0;
    assign fifo_intf_726.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_726;
    csv_file_dump cstatus_csv_dumper_726;
    df_fifo_monitor fifo_monitor_726;
    df_fifo_intf fifo_intf_727(clock,reset);
    assign fifo_intf_727.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_35_U.if_empty_n;
    assign fifo_intf_727.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_35_U.if_full_n;
    assign fifo_intf_727.fifo_rd_block = 0;
    assign fifo_intf_727.fifo_wr_block = 0;
    assign fifo_intf_727.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_727;
    csv_file_dump cstatus_csv_dumper_727;
    df_fifo_monitor fifo_monitor_727;
    df_fifo_intf fifo_intf_728(clock,reset);
    assign fifo_intf_728.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_35_U.if_empty_n;
    assign fifo_intf_728.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_35_U.if_full_n;
    assign fifo_intf_728.fifo_rd_block = 0;
    assign fifo_intf_728.fifo_wr_block = 0;
    assign fifo_intf_728.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_728;
    csv_file_dump cstatus_csv_dumper_728;
    df_fifo_monitor fifo_monitor_728;
    df_fifo_intf fifo_intf_729(clock,reset);
    assign fifo_intf_729.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_35_U.if_empty_n;
    assign fifo_intf_729.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_35_U.if_full_n;
    assign fifo_intf_729.fifo_rd_block = 0;
    assign fifo_intf_729.fifo_wr_block = 0;
    assign fifo_intf_729.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_729;
    csv_file_dump cstatus_csv_dumper_729;
    df_fifo_monitor fifo_monitor_729;
    df_fifo_intf fifo_intf_730(clock,reset);
    assign fifo_intf_730.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_35_U.if_empty_n;
    assign fifo_intf_730.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_35_U.if_full_n;
    assign fifo_intf_730.fifo_rd_block = 0;
    assign fifo_intf_730.fifo_wr_block = 0;
    assign fifo_intf_730.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_730;
    csv_file_dump cstatus_csv_dumper_730;
    df_fifo_monitor fifo_monitor_730;
    df_fifo_intf fifo_intf_731(clock,reset);
    assign fifo_intf_731.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_35_U.if_empty_n;
    assign fifo_intf_731.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_35_U.if_full_n;
    assign fifo_intf_731.fifo_rd_block = 0;
    assign fifo_intf_731.fifo_wr_block = 0;
    assign fifo_intf_731.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_731;
    csv_file_dump cstatus_csv_dumper_731;
    df_fifo_monitor fifo_monitor_731;
    df_fifo_intf fifo_intf_732(clock,reset);
    assign fifo_intf_732.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_35_U.if_empty_n;
    assign fifo_intf_732.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_35_U.if_full_n;
    assign fifo_intf_732.fifo_rd_block = 0;
    assign fifo_intf_732.fifo_wr_block = 0;
    assign fifo_intf_732.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_732;
    csv_file_dump cstatus_csv_dumper_732;
    df_fifo_monitor fifo_monitor_732;
    df_fifo_intf fifo_intf_733(clock,reset);
    assign fifo_intf_733.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_35_U.if_empty_n;
    assign fifo_intf_733.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_35_U.if_full_n;
    assign fifo_intf_733.fifo_rd_block = 0;
    assign fifo_intf_733.fifo_wr_block = 0;
    assign fifo_intf_733.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_733;
    csv_file_dump cstatus_csv_dumper_733;
    df_fifo_monitor fifo_monitor_733;
    df_fifo_intf fifo_intf_734(clock,reset);
    assign fifo_intf_734.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_35_U.if_empty_n;
    assign fifo_intf_734.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_35_U.if_full_n;
    assign fifo_intf_734.fifo_rd_block = 0;
    assign fifo_intf_734.fifo_wr_block = 0;
    assign fifo_intf_734.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_734;
    csv_file_dump cstatus_csv_dumper_734;
    df_fifo_monitor fifo_monitor_734;
    df_fifo_intf fifo_intf_735(clock,reset);
    assign fifo_intf_735.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_35_U.if_empty_n;
    assign fifo_intf_735.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_35_U.if_full_n;
    assign fifo_intf_735.fifo_rd_block = 0;
    assign fifo_intf_735.fifo_wr_block = 0;
    assign fifo_intf_735.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_735;
    csv_file_dump cstatus_csv_dumper_735;
    df_fifo_monitor fifo_monitor_735;
    df_fifo_intf fifo_intf_736(clock,reset);
    assign fifo_intf_736.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_35_U.if_empty_n;
    assign fifo_intf_736.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_35_U.if_full_n;
    assign fifo_intf_736.fifo_rd_block = 0;
    assign fifo_intf_736.fifo_wr_block = 0;
    assign fifo_intf_736.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_736;
    csv_file_dump cstatus_csv_dumper_736;
    df_fifo_monitor fifo_monitor_736;
    df_fifo_intf fifo_intf_737(clock,reset);
    assign fifo_intf_737.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_35_U.if_empty_n;
    assign fifo_intf_737.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_35_U.if_full_n;
    assign fifo_intf_737.fifo_rd_block = 0;
    assign fifo_intf_737.fifo_wr_block = 0;
    assign fifo_intf_737.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_737;
    csv_file_dump cstatus_csv_dumper_737;
    df_fifo_monitor fifo_monitor_737;
    df_fifo_intf fifo_intf_738(clock,reset);
    assign fifo_intf_738.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_35_U.if_empty_n;
    assign fifo_intf_738.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_35_U.if_full_n;
    assign fifo_intf_738.fifo_rd_block = 0;
    assign fifo_intf_738.fifo_wr_block = 0;
    assign fifo_intf_738.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_738;
    csv_file_dump cstatus_csv_dumper_738;
    df_fifo_monitor fifo_monitor_738;
    df_fifo_intf fifo_intf_739(clock,reset);
    assign fifo_intf_739.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_35_U.if_empty_n;
    assign fifo_intf_739.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_35_U.if_full_n;
    assign fifo_intf_739.fifo_rd_block = 0;
    assign fifo_intf_739.fifo_wr_block = 0;
    assign fifo_intf_739.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_739;
    csv_file_dump cstatus_csv_dumper_739;
    df_fifo_monitor fifo_monitor_739;
    df_fifo_intf fifo_intf_740(clock,reset);
    assign fifo_intf_740.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_35_U.if_empty_n;
    assign fifo_intf_740.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_35_U.if_full_n;
    assign fifo_intf_740.fifo_rd_block = 0;
    assign fifo_intf_740.fifo_wr_block = 0;
    assign fifo_intf_740.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_740;
    csv_file_dump cstatus_csv_dumper_740;
    df_fifo_monitor fifo_monitor_740;
    df_fifo_intf fifo_intf_741(clock,reset);
    assign fifo_intf_741.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_35_U.if_empty_n;
    assign fifo_intf_741.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_35_U.if_full_n;
    assign fifo_intf_741.fifo_rd_block = 0;
    assign fifo_intf_741.fifo_wr_block = 0;
    assign fifo_intf_741.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_741;
    csv_file_dump cstatus_csv_dumper_741;
    df_fifo_monitor fifo_monitor_741;
    df_fifo_intf fifo_intf_742(clock,reset);
    assign fifo_intf_742.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_35_U.if_empty_n;
    assign fifo_intf_742.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_35_U.if_full_n;
    assign fifo_intf_742.fifo_rd_block = 0;
    assign fifo_intf_742.fifo_wr_block = 0;
    assign fifo_intf_742.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_742;
    csv_file_dump cstatus_csv_dumper_742;
    df_fifo_monitor fifo_monitor_742;
    df_fifo_intf fifo_intf_743(clock,reset);
    assign fifo_intf_743.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_35_U.if_empty_n;
    assign fifo_intf_743.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_35_U.if_full_n;
    assign fifo_intf_743.fifo_rd_block = 0;
    assign fifo_intf_743.fifo_wr_block = 0;
    assign fifo_intf_743.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_743;
    csv_file_dump cstatus_csv_dumper_743;
    df_fifo_monitor fifo_monitor_743;
    df_fifo_intf fifo_intf_744(clock,reset);
    assign fifo_intf_744.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_35_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_35_U.if_empty_n;
    assign fifo_intf_744.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_35_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_35_U.if_full_n;
    assign fifo_intf_744.fifo_rd_block = 0;
    assign fifo_intf_744.fifo_wr_block = 0;
    assign fifo_intf_744.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_744;
    csv_file_dump cstatus_csv_dumper_744;
    df_fifo_monitor fifo_monitor_744;
    df_fifo_intf fifo_intf_745(clock,reset);
    assign fifo_intf_745.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_36_U.if_empty_n;
    assign fifo_intf_745.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_36_U.if_full_n;
    assign fifo_intf_745.fifo_rd_block = 0;
    assign fifo_intf_745.fifo_wr_block = 0;
    assign fifo_intf_745.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_745;
    csv_file_dump cstatus_csv_dumper_745;
    df_fifo_monitor fifo_monitor_745;
    df_fifo_intf fifo_intf_746(clock,reset);
    assign fifo_intf_746.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_36_U.if_empty_n;
    assign fifo_intf_746.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_36_U.if_full_n;
    assign fifo_intf_746.fifo_rd_block = 0;
    assign fifo_intf_746.fifo_wr_block = 0;
    assign fifo_intf_746.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_746;
    csv_file_dump cstatus_csv_dumper_746;
    df_fifo_monitor fifo_monitor_746;
    df_fifo_intf fifo_intf_747(clock,reset);
    assign fifo_intf_747.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_36_U.if_empty_n;
    assign fifo_intf_747.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_36_U.if_full_n;
    assign fifo_intf_747.fifo_rd_block = 0;
    assign fifo_intf_747.fifo_wr_block = 0;
    assign fifo_intf_747.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_747;
    csv_file_dump cstatus_csv_dumper_747;
    df_fifo_monitor fifo_monitor_747;
    df_fifo_intf fifo_intf_748(clock,reset);
    assign fifo_intf_748.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_36_U.if_empty_n;
    assign fifo_intf_748.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_36_U.if_full_n;
    assign fifo_intf_748.fifo_rd_block = 0;
    assign fifo_intf_748.fifo_wr_block = 0;
    assign fifo_intf_748.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_748;
    csv_file_dump cstatus_csv_dumper_748;
    df_fifo_monitor fifo_monitor_748;
    df_fifo_intf fifo_intf_749(clock,reset);
    assign fifo_intf_749.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_36_U.if_empty_n;
    assign fifo_intf_749.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_36_U.if_full_n;
    assign fifo_intf_749.fifo_rd_block = 0;
    assign fifo_intf_749.fifo_wr_block = 0;
    assign fifo_intf_749.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_749;
    csv_file_dump cstatus_csv_dumper_749;
    df_fifo_monitor fifo_monitor_749;
    df_fifo_intf fifo_intf_750(clock,reset);
    assign fifo_intf_750.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_36_U.if_empty_n;
    assign fifo_intf_750.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_36_U.if_full_n;
    assign fifo_intf_750.fifo_rd_block = 0;
    assign fifo_intf_750.fifo_wr_block = 0;
    assign fifo_intf_750.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_750;
    csv_file_dump cstatus_csv_dumper_750;
    df_fifo_monitor fifo_monitor_750;
    df_fifo_intf fifo_intf_751(clock,reset);
    assign fifo_intf_751.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_36_U.if_empty_n;
    assign fifo_intf_751.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_36_U.if_full_n;
    assign fifo_intf_751.fifo_rd_block = 0;
    assign fifo_intf_751.fifo_wr_block = 0;
    assign fifo_intf_751.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_751;
    csv_file_dump cstatus_csv_dumper_751;
    df_fifo_monitor fifo_monitor_751;
    df_fifo_intf fifo_intf_752(clock,reset);
    assign fifo_intf_752.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_36_U.if_empty_n;
    assign fifo_intf_752.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_36_U.if_full_n;
    assign fifo_intf_752.fifo_rd_block = 0;
    assign fifo_intf_752.fifo_wr_block = 0;
    assign fifo_intf_752.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_752;
    csv_file_dump cstatus_csv_dumper_752;
    df_fifo_monitor fifo_monitor_752;
    df_fifo_intf fifo_intf_753(clock,reset);
    assign fifo_intf_753.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_36_U.if_empty_n;
    assign fifo_intf_753.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_36_U.if_full_n;
    assign fifo_intf_753.fifo_rd_block = 0;
    assign fifo_intf_753.fifo_wr_block = 0;
    assign fifo_intf_753.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_753;
    csv_file_dump cstatus_csv_dumper_753;
    df_fifo_monitor fifo_monitor_753;
    df_fifo_intf fifo_intf_754(clock,reset);
    assign fifo_intf_754.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_36_U.if_empty_n;
    assign fifo_intf_754.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_36_U.if_full_n;
    assign fifo_intf_754.fifo_rd_block = 0;
    assign fifo_intf_754.fifo_wr_block = 0;
    assign fifo_intf_754.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_754;
    csv_file_dump cstatus_csv_dumper_754;
    df_fifo_monitor fifo_monitor_754;
    df_fifo_intf fifo_intf_755(clock,reset);
    assign fifo_intf_755.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_36_U.if_empty_n;
    assign fifo_intf_755.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_36_U.if_full_n;
    assign fifo_intf_755.fifo_rd_block = 0;
    assign fifo_intf_755.fifo_wr_block = 0;
    assign fifo_intf_755.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_755;
    csv_file_dump cstatus_csv_dumper_755;
    df_fifo_monitor fifo_monitor_755;
    df_fifo_intf fifo_intf_756(clock,reset);
    assign fifo_intf_756.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_36_U.if_empty_n;
    assign fifo_intf_756.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_36_U.if_full_n;
    assign fifo_intf_756.fifo_rd_block = 0;
    assign fifo_intf_756.fifo_wr_block = 0;
    assign fifo_intf_756.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_756;
    csv_file_dump cstatus_csv_dumper_756;
    df_fifo_monitor fifo_monitor_756;
    df_fifo_intf fifo_intf_757(clock,reset);
    assign fifo_intf_757.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_36_U.if_empty_n;
    assign fifo_intf_757.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_36_U.if_full_n;
    assign fifo_intf_757.fifo_rd_block = 0;
    assign fifo_intf_757.fifo_wr_block = 0;
    assign fifo_intf_757.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_757;
    csv_file_dump cstatus_csv_dumper_757;
    df_fifo_monitor fifo_monitor_757;
    df_fifo_intf fifo_intf_758(clock,reset);
    assign fifo_intf_758.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_36_U.if_empty_n;
    assign fifo_intf_758.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_36_U.if_full_n;
    assign fifo_intf_758.fifo_rd_block = 0;
    assign fifo_intf_758.fifo_wr_block = 0;
    assign fifo_intf_758.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_758;
    csv_file_dump cstatus_csv_dumper_758;
    df_fifo_monitor fifo_monitor_758;
    df_fifo_intf fifo_intf_759(clock,reset);
    assign fifo_intf_759.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_36_U.if_empty_n;
    assign fifo_intf_759.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_36_U.if_full_n;
    assign fifo_intf_759.fifo_rd_block = 0;
    assign fifo_intf_759.fifo_wr_block = 0;
    assign fifo_intf_759.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_759;
    csv_file_dump cstatus_csv_dumper_759;
    df_fifo_monitor fifo_monitor_759;
    df_fifo_intf fifo_intf_760(clock,reset);
    assign fifo_intf_760.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_36_U.if_empty_n;
    assign fifo_intf_760.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_36_U.if_full_n;
    assign fifo_intf_760.fifo_rd_block = 0;
    assign fifo_intf_760.fifo_wr_block = 0;
    assign fifo_intf_760.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_760;
    csv_file_dump cstatus_csv_dumper_760;
    df_fifo_monitor fifo_monitor_760;
    df_fifo_intf fifo_intf_761(clock,reset);
    assign fifo_intf_761.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_36_U.if_empty_n;
    assign fifo_intf_761.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_36_U.if_full_n;
    assign fifo_intf_761.fifo_rd_block = 0;
    assign fifo_intf_761.fifo_wr_block = 0;
    assign fifo_intf_761.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_761;
    csv_file_dump cstatus_csv_dumper_761;
    df_fifo_monitor fifo_monitor_761;
    df_fifo_intf fifo_intf_762(clock,reset);
    assign fifo_intf_762.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_36_U.if_empty_n;
    assign fifo_intf_762.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_36_U.if_full_n;
    assign fifo_intf_762.fifo_rd_block = 0;
    assign fifo_intf_762.fifo_wr_block = 0;
    assign fifo_intf_762.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_762;
    csv_file_dump cstatus_csv_dumper_762;
    df_fifo_monitor fifo_monitor_762;
    df_fifo_intf fifo_intf_763(clock,reset);
    assign fifo_intf_763.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_36_U.if_empty_n;
    assign fifo_intf_763.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_36_U.if_full_n;
    assign fifo_intf_763.fifo_rd_block = 0;
    assign fifo_intf_763.fifo_wr_block = 0;
    assign fifo_intf_763.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_763;
    csv_file_dump cstatus_csv_dumper_763;
    df_fifo_monitor fifo_monitor_763;
    df_fifo_intf fifo_intf_764(clock,reset);
    assign fifo_intf_764.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_36_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_36_U.if_empty_n;
    assign fifo_intf_764.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_36_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_36_U.if_full_n;
    assign fifo_intf_764.fifo_rd_block = 0;
    assign fifo_intf_764.fifo_wr_block = 0;
    assign fifo_intf_764.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_764;
    csv_file_dump cstatus_csv_dumper_764;
    df_fifo_monitor fifo_monitor_764;
    df_fifo_intf fifo_intf_765(clock,reset);
    assign fifo_intf_765.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_37_U.if_empty_n;
    assign fifo_intf_765.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_37_U.if_full_n;
    assign fifo_intf_765.fifo_rd_block = 0;
    assign fifo_intf_765.fifo_wr_block = 0;
    assign fifo_intf_765.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_765;
    csv_file_dump cstatus_csv_dumper_765;
    df_fifo_monitor fifo_monitor_765;
    df_fifo_intf fifo_intf_766(clock,reset);
    assign fifo_intf_766.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_37_U.if_empty_n;
    assign fifo_intf_766.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_37_U.if_full_n;
    assign fifo_intf_766.fifo_rd_block = 0;
    assign fifo_intf_766.fifo_wr_block = 0;
    assign fifo_intf_766.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_766;
    csv_file_dump cstatus_csv_dumper_766;
    df_fifo_monitor fifo_monitor_766;
    df_fifo_intf fifo_intf_767(clock,reset);
    assign fifo_intf_767.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_37_U.if_empty_n;
    assign fifo_intf_767.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_37_U.if_full_n;
    assign fifo_intf_767.fifo_rd_block = 0;
    assign fifo_intf_767.fifo_wr_block = 0;
    assign fifo_intf_767.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_767;
    csv_file_dump cstatus_csv_dumper_767;
    df_fifo_monitor fifo_monitor_767;
    df_fifo_intf fifo_intf_768(clock,reset);
    assign fifo_intf_768.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_37_U.if_empty_n;
    assign fifo_intf_768.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_37_U.if_full_n;
    assign fifo_intf_768.fifo_rd_block = 0;
    assign fifo_intf_768.fifo_wr_block = 0;
    assign fifo_intf_768.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_768;
    csv_file_dump cstatus_csv_dumper_768;
    df_fifo_monitor fifo_monitor_768;
    df_fifo_intf fifo_intf_769(clock,reset);
    assign fifo_intf_769.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_37_U.if_empty_n;
    assign fifo_intf_769.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_37_U.if_full_n;
    assign fifo_intf_769.fifo_rd_block = 0;
    assign fifo_intf_769.fifo_wr_block = 0;
    assign fifo_intf_769.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_769;
    csv_file_dump cstatus_csv_dumper_769;
    df_fifo_monitor fifo_monitor_769;
    df_fifo_intf fifo_intf_770(clock,reset);
    assign fifo_intf_770.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_37_U.if_empty_n;
    assign fifo_intf_770.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_37_U.if_full_n;
    assign fifo_intf_770.fifo_rd_block = 0;
    assign fifo_intf_770.fifo_wr_block = 0;
    assign fifo_intf_770.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_770;
    csv_file_dump cstatus_csv_dumper_770;
    df_fifo_monitor fifo_monitor_770;
    df_fifo_intf fifo_intf_771(clock,reset);
    assign fifo_intf_771.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_37_U.if_empty_n;
    assign fifo_intf_771.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_37_U.if_full_n;
    assign fifo_intf_771.fifo_rd_block = 0;
    assign fifo_intf_771.fifo_wr_block = 0;
    assign fifo_intf_771.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_771;
    csv_file_dump cstatus_csv_dumper_771;
    df_fifo_monitor fifo_monitor_771;
    df_fifo_intf fifo_intf_772(clock,reset);
    assign fifo_intf_772.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_37_U.if_empty_n;
    assign fifo_intf_772.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_37_U.if_full_n;
    assign fifo_intf_772.fifo_rd_block = 0;
    assign fifo_intf_772.fifo_wr_block = 0;
    assign fifo_intf_772.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_772;
    csv_file_dump cstatus_csv_dumper_772;
    df_fifo_monitor fifo_monitor_772;
    df_fifo_intf fifo_intf_773(clock,reset);
    assign fifo_intf_773.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_37_U.if_empty_n;
    assign fifo_intf_773.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_37_U.if_full_n;
    assign fifo_intf_773.fifo_rd_block = 0;
    assign fifo_intf_773.fifo_wr_block = 0;
    assign fifo_intf_773.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_773;
    csv_file_dump cstatus_csv_dumper_773;
    df_fifo_monitor fifo_monitor_773;
    df_fifo_intf fifo_intf_774(clock,reset);
    assign fifo_intf_774.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_37_U.if_empty_n;
    assign fifo_intf_774.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_37_U.if_full_n;
    assign fifo_intf_774.fifo_rd_block = 0;
    assign fifo_intf_774.fifo_wr_block = 0;
    assign fifo_intf_774.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_774;
    csv_file_dump cstatus_csv_dumper_774;
    df_fifo_monitor fifo_monitor_774;
    df_fifo_intf fifo_intf_775(clock,reset);
    assign fifo_intf_775.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_37_U.if_empty_n;
    assign fifo_intf_775.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_37_U.if_full_n;
    assign fifo_intf_775.fifo_rd_block = 0;
    assign fifo_intf_775.fifo_wr_block = 0;
    assign fifo_intf_775.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_775;
    csv_file_dump cstatus_csv_dumper_775;
    df_fifo_monitor fifo_monitor_775;
    df_fifo_intf fifo_intf_776(clock,reset);
    assign fifo_intf_776.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_37_U.if_empty_n;
    assign fifo_intf_776.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_37_U.if_full_n;
    assign fifo_intf_776.fifo_rd_block = 0;
    assign fifo_intf_776.fifo_wr_block = 0;
    assign fifo_intf_776.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_776;
    csv_file_dump cstatus_csv_dumper_776;
    df_fifo_monitor fifo_monitor_776;
    df_fifo_intf fifo_intf_777(clock,reset);
    assign fifo_intf_777.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_37_U.if_empty_n;
    assign fifo_intf_777.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_37_U.if_full_n;
    assign fifo_intf_777.fifo_rd_block = 0;
    assign fifo_intf_777.fifo_wr_block = 0;
    assign fifo_intf_777.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_777;
    csv_file_dump cstatus_csv_dumper_777;
    df_fifo_monitor fifo_monitor_777;
    df_fifo_intf fifo_intf_778(clock,reset);
    assign fifo_intf_778.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_37_U.if_empty_n;
    assign fifo_intf_778.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_37_U.if_full_n;
    assign fifo_intf_778.fifo_rd_block = 0;
    assign fifo_intf_778.fifo_wr_block = 0;
    assign fifo_intf_778.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_778;
    csv_file_dump cstatus_csv_dumper_778;
    df_fifo_monitor fifo_monitor_778;
    df_fifo_intf fifo_intf_779(clock,reset);
    assign fifo_intf_779.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_37_U.if_empty_n;
    assign fifo_intf_779.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_37_U.if_full_n;
    assign fifo_intf_779.fifo_rd_block = 0;
    assign fifo_intf_779.fifo_wr_block = 0;
    assign fifo_intf_779.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_779;
    csv_file_dump cstatus_csv_dumper_779;
    df_fifo_monitor fifo_monitor_779;
    df_fifo_intf fifo_intf_780(clock,reset);
    assign fifo_intf_780.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_37_U.if_empty_n;
    assign fifo_intf_780.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_37_U.if_full_n;
    assign fifo_intf_780.fifo_rd_block = 0;
    assign fifo_intf_780.fifo_wr_block = 0;
    assign fifo_intf_780.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_780;
    csv_file_dump cstatus_csv_dumper_780;
    df_fifo_monitor fifo_monitor_780;
    df_fifo_intf fifo_intf_781(clock,reset);
    assign fifo_intf_781.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_37_U.if_empty_n;
    assign fifo_intf_781.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_37_U.if_full_n;
    assign fifo_intf_781.fifo_rd_block = 0;
    assign fifo_intf_781.fifo_wr_block = 0;
    assign fifo_intf_781.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_781;
    csv_file_dump cstatus_csv_dumper_781;
    df_fifo_monitor fifo_monitor_781;
    df_fifo_intf fifo_intf_782(clock,reset);
    assign fifo_intf_782.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_37_U.if_empty_n;
    assign fifo_intf_782.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_37_U.if_full_n;
    assign fifo_intf_782.fifo_rd_block = 0;
    assign fifo_intf_782.fifo_wr_block = 0;
    assign fifo_intf_782.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_782;
    csv_file_dump cstatus_csv_dumper_782;
    df_fifo_monitor fifo_monitor_782;
    df_fifo_intf fifo_intf_783(clock,reset);
    assign fifo_intf_783.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_37_U.if_empty_n;
    assign fifo_intf_783.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_37_U.if_full_n;
    assign fifo_intf_783.fifo_rd_block = 0;
    assign fifo_intf_783.fifo_wr_block = 0;
    assign fifo_intf_783.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_783;
    csv_file_dump cstatus_csv_dumper_783;
    df_fifo_monitor fifo_monitor_783;
    df_fifo_intf fifo_intf_784(clock,reset);
    assign fifo_intf_784.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_37_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_37_U.if_empty_n;
    assign fifo_intf_784.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_37_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_37_U.if_full_n;
    assign fifo_intf_784.fifo_rd_block = 0;
    assign fifo_intf_784.fifo_wr_block = 0;
    assign fifo_intf_784.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_784;
    csv_file_dump cstatus_csv_dumper_784;
    df_fifo_monitor fifo_monitor_784;
    df_fifo_intf fifo_intf_785(clock,reset);
    assign fifo_intf_785.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_38_U.if_empty_n;
    assign fifo_intf_785.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_38_U.if_full_n;
    assign fifo_intf_785.fifo_rd_block = 0;
    assign fifo_intf_785.fifo_wr_block = 0;
    assign fifo_intf_785.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_785;
    csv_file_dump cstatus_csv_dumper_785;
    df_fifo_monitor fifo_monitor_785;
    df_fifo_intf fifo_intf_786(clock,reset);
    assign fifo_intf_786.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_38_U.if_empty_n;
    assign fifo_intf_786.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_38_U.if_full_n;
    assign fifo_intf_786.fifo_rd_block = 0;
    assign fifo_intf_786.fifo_wr_block = 0;
    assign fifo_intf_786.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_786;
    csv_file_dump cstatus_csv_dumper_786;
    df_fifo_monitor fifo_monitor_786;
    df_fifo_intf fifo_intf_787(clock,reset);
    assign fifo_intf_787.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_38_U.if_empty_n;
    assign fifo_intf_787.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_38_U.if_full_n;
    assign fifo_intf_787.fifo_rd_block = 0;
    assign fifo_intf_787.fifo_wr_block = 0;
    assign fifo_intf_787.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_787;
    csv_file_dump cstatus_csv_dumper_787;
    df_fifo_monitor fifo_monitor_787;
    df_fifo_intf fifo_intf_788(clock,reset);
    assign fifo_intf_788.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_38_U.if_empty_n;
    assign fifo_intf_788.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_38_U.if_full_n;
    assign fifo_intf_788.fifo_rd_block = 0;
    assign fifo_intf_788.fifo_wr_block = 0;
    assign fifo_intf_788.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_788;
    csv_file_dump cstatus_csv_dumper_788;
    df_fifo_monitor fifo_monitor_788;
    df_fifo_intf fifo_intf_789(clock,reset);
    assign fifo_intf_789.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_38_U.if_empty_n;
    assign fifo_intf_789.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_38_U.if_full_n;
    assign fifo_intf_789.fifo_rd_block = 0;
    assign fifo_intf_789.fifo_wr_block = 0;
    assign fifo_intf_789.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_789;
    csv_file_dump cstatus_csv_dumper_789;
    df_fifo_monitor fifo_monitor_789;
    df_fifo_intf fifo_intf_790(clock,reset);
    assign fifo_intf_790.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_38_U.if_empty_n;
    assign fifo_intf_790.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_38_U.if_full_n;
    assign fifo_intf_790.fifo_rd_block = 0;
    assign fifo_intf_790.fifo_wr_block = 0;
    assign fifo_intf_790.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_790;
    csv_file_dump cstatus_csv_dumper_790;
    df_fifo_monitor fifo_monitor_790;
    df_fifo_intf fifo_intf_791(clock,reset);
    assign fifo_intf_791.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_38_U.if_empty_n;
    assign fifo_intf_791.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_38_U.if_full_n;
    assign fifo_intf_791.fifo_rd_block = 0;
    assign fifo_intf_791.fifo_wr_block = 0;
    assign fifo_intf_791.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_791;
    csv_file_dump cstatus_csv_dumper_791;
    df_fifo_monitor fifo_monitor_791;
    df_fifo_intf fifo_intf_792(clock,reset);
    assign fifo_intf_792.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_38_U.if_empty_n;
    assign fifo_intf_792.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_38_U.if_full_n;
    assign fifo_intf_792.fifo_rd_block = 0;
    assign fifo_intf_792.fifo_wr_block = 0;
    assign fifo_intf_792.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_792;
    csv_file_dump cstatus_csv_dumper_792;
    df_fifo_monitor fifo_monitor_792;
    df_fifo_intf fifo_intf_793(clock,reset);
    assign fifo_intf_793.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_38_U.if_empty_n;
    assign fifo_intf_793.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_38_U.if_full_n;
    assign fifo_intf_793.fifo_rd_block = 0;
    assign fifo_intf_793.fifo_wr_block = 0;
    assign fifo_intf_793.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_793;
    csv_file_dump cstatus_csv_dumper_793;
    df_fifo_monitor fifo_monitor_793;
    df_fifo_intf fifo_intf_794(clock,reset);
    assign fifo_intf_794.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_38_U.if_empty_n;
    assign fifo_intf_794.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_38_U.if_full_n;
    assign fifo_intf_794.fifo_rd_block = 0;
    assign fifo_intf_794.fifo_wr_block = 0;
    assign fifo_intf_794.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_794;
    csv_file_dump cstatus_csv_dumper_794;
    df_fifo_monitor fifo_monitor_794;
    df_fifo_intf fifo_intf_795(clock,reset);
    assign fifo_intf_795.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_38_U.if_empty_n;
    assign fifo_intf_795.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_38_U.if_full_n;
    assign fifo_intf_795.fifo_rd_block = 0;
    assign fifo_intf_795.fifo_wr_block = 0;
    assign fifo_intf_795.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_795;
    csv_file_dump cstatus_csv_dumper_795;
    df_fifo_monitor fifo_monitor_795;
    df_fifo_intf fifo_intf_796(clock,reset);
    assign fifo_intf_796.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_38_U.if_empty_n;
    assign fifo_intf_796.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_38_U.if_full_n;
    assign fifo_intf_796.fifo_rd_block = 0;
    assign fifo_intf_796.fifo_wr_block = 0;
    assign fifo_intf_796.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_796;
    csv_file_dump cstatus_csv_dumper_796;
    df_fifo_monitor fifo_monitor_796;
    df_fifo_intf fifo_intf_797(clock,reset);
    assign fifo_intf_797.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_38_U.if_empty_n;
    assign fifo_intf_797.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_38_U.if_full_n;
    assign fifo_intf_797.fifo_rd_block = 0;
    assign fifo_intf_797.fifo_wr_block = 0;
    assign fifo_intf_797.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_797;
    csv_file_dump cstatus_csv_dumper_797;
    df_fifo_monitor fifo_monitor_797;
    df_fifo_intf fifo_intf_798(clock,reset);
    assign fifo_intf_798.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_38_U.if_empty_n;
    assign fifo_intf_798.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_38_U.if_full_n;
    assign fifo_intf_798.fifo_rd_block = 0;
    assign fifo_intf_798.fifo_wr_block = 0;
    assign fifo_intf_798.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_798;
    csv_file_dump cstatus_csv_dumper_798;
    df_fifo_monitor fifo_monitor_798;
    df_fifo_intf fifo_intf_799(clock,reset);
    assign fifo_intf_799.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_38_U.if_empty_n;
    assign fifo_intf_799.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_38_U.if_full_n;
    assign fifo_intf_799.fifo_rd_block = 0;
    assign fifo_intf_799.fifo_wr_block = 0;
    assign fifo_intf_799.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_799;
    csv_file_dump cstatus_csv_dumper_799;
    df_fifo_monitor fifo_monitor_799;
    df_fifo_intf fifo_intf_800(clock,reset);
    assign fifo_intf_800.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_38_U.if_empty_n;
    assign fifo_intf_800.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_38_U.if_full_n;
    assign fifo_intf_800.fifo_rd_block = 0;
    assign fifo_intf_800.fifo_wr_block = 0;
    assign fifo_intf_800.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_800;
    csv_file_dump cstatus_csv_dumper_800;
    df_fifo_monitor fifo_monitor_800;
    df_fifo_intf fifo_intf_801(clock,reset);
    assign fifo_intf_801.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_38_U.if_empty_n;
    assign fifo_intf_801.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_38_U.if_full_n;
    assign fifo_intf_801.fifo_rd_block = 0;
    assign fifo_intf_801.fifo_wr_block = 0;
    assign fifo_intf_801.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_801;
    csv_file_dump cstatus_csv_dumper_801;
    df_fifo_monitor fifo_monitor_801;
    df_fifo_intf fifo_intf_802(clock,reset);
    assign fifo_intf_802.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_38_U.if_empty_n;
    assign fifo_intf_802.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_38_U.if_full_n;
    assign fifo_intf_802.fifo_rd_block = 0;
    assign fifo_intf_802.fifo_wr_block = 0;
    assign fifo_intf_802.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_802;
    csv_file_dump cstatus_csv_dumper_802;
    df_fifo_monitor fifo_monitor_802;
    df_fifo_intf fifo_intf_803(clock,reset);
    assign fifo_intf_803.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_38_U.if_empty_n;
    assign fifo_intf_803.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_38_U.if_full_n;
    assign fifo_intf_803.fifo_rd_block = 0;
    assign fifo_intf_803.fifo_wr_block = 0;
    assign fifo_intf_803.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_803;
    csv_file_dump cstatus_csv_dumper_803;
    df_fifo_monitor fifo_monitor_803;
    df_fifo_intf fifo_intf_804(clock,reset);
    assign fifo_intf_804.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_38_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_38_U.if_empty_n;
    assign fifo_intf_804.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_38_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_38_U.if_full_n;
    assign fifo_intf_804.fifo_rd_block = 0;
    assign fifo_intf_804.fifo_wr_block = 0;
    assign fifo_intf_804.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_804;
    csv_file_dump cstatus_csv_dumper_804;
    df_fifo_monitor fifo_monitor_804;
    df_fifo_intf fifo_intf_805(clock,reset);
    assign fifo_intf_805.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_39_U.if_empty_n;
    assign fifo_intf_805.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_0_39_U.if_full_n;
    assign fifo_intf_805.fifo_rd_block = 0;
    assign fifo_intf_805.fifo_wr_block = 0;
    assign fifo_intf_805.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_805;
    csv_file_dump cstatus_csv_dumper_805;
    df_fifo_monitor fifo_monitor_805;
    df_fifo_intf fifo_intf_806(clock,reset);
    assign fifo_intf_806.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_39_U.if_empty_n;
    assign fifo_intf_806.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_1_39_U.if_full_n;
    assign fifo_intf_806.fifo_rd_block = 0;
    assign fifo_intf_806.fifo_wr_block = 0;
    assign fifo_intf_806.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_806;
    csv_file_dump cstatus_csv_dumper_806;
    df_fifo_monitor fifo_monitor_806;
    df_fifo_intf fifo_intf_807(clock,reset);
    assign fifo_intf_807.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_39_U.if_empty_n;
    assign fifo_intf_807.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_2_39_U.if_full_n;
    assign fifo_intf_807.fifo_rd_block = 0;
    assign fifo_intf_807.fifo_wr_block = 0;
    assign fifo_intf_807.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_807;
    csv_file_dump cstatus_csv_dumper_807;
    df_fifo_monitor fifo_monitor_807;
    df_fifo_intf fifo_intf_808(clock,reset);
    assign fifo_intf_808.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_39_U.if_empty_n;
    assign fifo_intf_808.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_3_39_U.if_full_n;
    assign fifo_intf_808.fifo_rd_block = 0;
    assign fifo_intf_808.fifo_wr_block = 0;
    assign fifo_intf_808.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_808;
    csv_file_dump cstatus_csv_dumper_808;
    df_fifo_monitor fifo_monitor_808;
    df_fifo_intf fifo_intf_809(clock,reset);
    assign fifo_intf_809.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_39_U.if_empty_n;
    assign fifo_intf_809.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_4_39_U.if_full_n;
    assign fifo_intf_809.fifo_rd_block = 0;
    assign fifo_intf_809.fifo_wr_block = 0;
    assign fifo_intf_809.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_809;
    csv_file_dump cstatus_csv_dumper_809;
    df_fifo_monitor fifo_monitor_809;
    df_fifo_intf fifo_intf_810(clock,reset);
    assign fifo_intf_810.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_39_U.if_empty_n;
    assign fifo_intf_810.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_5_39_U.if_full_n;
    assign fifo_intf_810.fifo_rd_block = 0;
    assign fifo_intf_810.fifo_wr_block = 0;
    assign fifo_intf_810.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_810;
    csv_file_dump cstatus_csv_dumper_810;
    df_fifo_monitor fifo_monitor_810;
    df_fifo_intf fifo_intf_811(clock,reset);
    assign fifo_intf_811.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_39_U.if_empty_n;
    assign fifo_intf_811.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_6_39_U.if_full_n;
    assign fifo_intf_811.fifo_rd_block = 0;
    assign fifo_intf_811.fifo_wr_block = 0;
    assign fifo_intf_811.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_811;
    csv_file_dump cstatus_csv_dumper_811;
    df_fifo_monitor fifo_monitor_811;
    df_fifo_intf fifo_intf_812(clock,reset);
    assign fifo_intf_812.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_39_U.if_empty_n;
    assign fifo_intf_812.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_7_39_U.if_full_n;
    assign fifo_intf_812.fifo_rd_block = 0;
    assign fifo_intf_812.fifo_wr_block = 0;
    assign fifo_intf_812.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_812;
    csv_file_dump cstatus_csv_dumper_812;
    df_fifo_monitor fifo_monitor_812;
    df_fifo_intf fifo_intf_813(clock,reset);
    assign fifo_intf_813.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_39_U.if_empty_n;
    assign fifo_intf_813.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_8_39_U.if_full_n;
    assign fifo_intf_813.fifo_rd_block = 0;
    assign fifo_intf_813.fifo_wr_block = 0;
    assign fifo_intf_813.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_813;
    csv_file_dump cstatus_csv_dumper_813;
    df_fifo_monitor fifo_monitor_813;
    df_fifo_intf fifo_intf_814(clock,reset);
    assign fifo_intf_814.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_39_U.if_empty_n;
    assign fifo_intf_814.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_9_39_U.if_full_n;
    assign fifo_intf_814.fifo_rd_block = 0;
    assign fifo_intf_814.fifo_wr_block = 0;
    assign fifo_intf_814.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_814;
    csv_file_dump cstatus_csv_dumper_814;
    df_fifo_monitor fifo_monitor_814;
    df_fifo_intf fifo_intf_815(clock,reset);
    assign fifo_intf_815.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_39_U.if_empty_n;
    assign fifo_intf_815.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_10_39_U.if_full_n;
    assign fifo_intf_815.fifo_rd_block = 0;
    assign fifo_intf_815.fifo_wr_block = 0;
    assign fifo_intf_815.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_815;
    csv_file_dump cstatus_csv_dumper_815;
    df_fifo_monitor fifo_monitor_815;
    df_fifo_intf fifo_intf_816(clock,reset);
    assign fifo_intf_816.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_39_U.if_empty_n;
    assign fifo_intf_816.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_11_39_U.if_full_n;
    assign fifo_intf_816.fifo_rd_block = 0;
    assign fifo_intf_816.fifo_wr_block = 0;
    assign fifo_intf_816.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_816;
    csv_file_dump cstatus_csv_dumper_816;
    df_fifo_monitor fifo_monitor_816;
    df_fifo_intf fifo_intf_817(clock,reset);
    assign fifo_intf_817.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_39_U.if_empty_n;
    assign fifo_intf_817.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_12_39_U.if_full_n;
    assign fifo_intf_817.fifo_rd_block = 0;
    assign fifo_intf_817.fifo_wr_block = 0;
    assign fifo_intf_817.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_817;
    csv_file_dump cstatus_csv_dumper_817;
    df_fifo_monitor fifo_monitor_817;
    df_fifo_intf fifo_intf_818(clock,reset);
    assign fifo_intf_818.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_39_U.if_empty_n;
    assign fifo_intf_818.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_13_39_U.if_full_n;
    assign fifo_intf_818.fifo_rd_block = 0;
    assign fifo_intf_818.fifo_wr_block = 0;
    assign fifo_intf_818.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_818;
    csv_file_dump cstatus_csv_dumper_818;
    df_fifo_monitor fifo_monitor_818;
    df_fifo_intf fifo_intf_819(clock,reset);
    assign fifo_intf_819.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_39_U.if_empty_n;
    assign fifo_intf_819.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_14_39_U.if_full_n;
    assign fifo_intf_819.fifo_rd_block = 0;
    assign fifo_intf_819.fifo_wr_block = 0;
    assign fifo_intf_819.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_819;
    csv_file_dump cstatus_csv_dumper_819;
    df_fifo_monitor fifo_monitor_819;
    df_fifo_intf fifo_intf_820(clock,reset);
    assign fifo_intf_820.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_39_U.if_empty_n;
    assign fifo_intf_820.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_15_39_U.if_full_n;
    assign fifo_intf_820.fifo_rd_block = 0;
    assign fifo_intf_820.fifo_wr_block = 0;
    assign fifo_intf_820.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_820;
    csv_file_dump cstatus_csv_dumper_820;
    df_fifo_monitor fifo_monitor_820;
    df_fifo_intf fifo_intf_821(clock,reset);
    assign fifo_intf_821.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_39_U.if_empty_n;
    assign fifo_intf_821.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_16_39_U.if_full_n;
    assign fifo_intf_821.fifo_rd_block = 0;
    assign fifo_intf_821.fifo_wr_block = 0;
    assign fifo_intf_821.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_821;
    csv_file_dump cstatus_csv_dumper_821;
    df_fifo_monitor fifo_monitor_821;
    df_fifo_intf fifo_intf_822(clock,reset);
    assign fifo_intf_822.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_39_U.if_empty_n;
    assign fifo_intf_822.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_17_39_U.if_full_n;
    assign fifo_intf_822.fifo_rd_block = 0;
    assign fifo_intf_822.fifo_wr_block = 0;
    assign fifo_intf_822.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_822;
    csv_file_dump cstatus_csv_dumper_822;
    df_fifo_monitor fifo_monitor_822;
    df_fifo_intf fifo_intf_823(clock,reset);
    assign fifo_intf_823.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_39_U.if_empty_n;
    assign fifo_intf_823.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_18_39_U.if_full_n;
    assign fifo_intf_823.fifo_rd_block = 0;
    assign fifo_intf_823.fifo_wr_block = 0;
    assign fifo_intf_823.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_823;
    csv_file_dump cstatus_csv_dumper_823;
    df_fifo_monitor fifo_monitor_823;
    df_fifo_intf fifo_intf_824(clock,reset);
    assign fifo_intf_824.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_39_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_39_U.if_empty_n;
    assign fifo_intf_824.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_39_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.qk_mul_19_39_U.if_full_n;
    assign fifo_intf_824.fifo_rd_block = 0;
    assign fifo_intf_824.fifo_wr_block = 0;
    assign fifo_intf_824.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_824;
    csv_file_dump cstatus_csv_dumper_824;
    df_fifo_monitor fifo_monitor_824;
    df_fifo_intf fifo_intf_825(clock,reset);
    assign fifo_intf_825.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_2_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_2_U.if_empty_n;
    assign fifo_intf_825.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_2_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_2_U.if_full_n;
    assign fifo_intf_825.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_0_blk_n);
    assign fifo_intf_825.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_0_blk_n);
    assign fifo_intf_825.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_825;
    csv_file_dump cstatus_csv_dumper_825;
    df_fifo_monitor fifo_monitor_825;
    df_fifo_intf fifo_intf_826(clock,reset);
    assign fifo_intf_826.rd_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_3_U.if_read & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_3_U.if_empty_n;
    assign fifo_intf_826.wr_en = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_3_U.if_write & AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matr_out_3_U.if_full_n;
    assign fifo_intf_826.fifo_rd_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_1_blk_n);
    assign fifo_intf_826.fifo_wr_block = ~(AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_1_blk_n);
    assign fifo_intf_826.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_826;
    csv_file_dump cstatus_csv_dumper_826;
    df_fifo_monitor fifo_monitor_826;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_myproject.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_myproject.ap_start == 1'b1 && AESL_inst_myproject.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_myproject.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end

logic region_1_idle;
logic [31:0] region_1_start_cnt;
logic [31:0] region_1_done_cnt;
assign region_1_idle = (region_1_start_cnt == region_1_done_cnt) && AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_start_cnt <= 32'h0;
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_start == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_ready == 1'b1)
        region_1_start_cnt <= region_1_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_done_cnt <= 32'h0;
    else if (AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_done == 1'b1 && AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_continue == 1'b1)
        region_1_done_cnt <= region_1_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.real_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_3_U0.d_query_0_3_blk_n;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_1_idle;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.real_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_2_U0.d_query_1_3_blk_n;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_1_idle;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_start;
    assign process_intf_3.pin_stall = 1'b0;
    assign process_intf_3.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_3_blk_n;
    assign process_intf_3.cin_stall = 1'b0;
    assign process_intf_3.cout_stall = 1'b0;
    assign process_intf_3.region_idle = region_1_idle;
    assign process_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_4.pin_stall = 1'b0;
    assign process_intf_4.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.data_prep_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_3_blk_n;
    assign process_intf_4.cin_stall = 1'b0;
    assign process_intf_4.cout_stall = 1'b0;
    assign process_intf_4.region_idle = region_1_idle;
    assign process_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.real_start;
    assign process_intf_5.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_query_0_3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.d_value_0_3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_3_blk_n;
    assign process_intf_5.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.k_proj_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.q_proj_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.v_proj_0_blk_n;
    assign process_intf_5.cin_stall = 1'b0;
    assign process_intf_5.cout_stall = 1'b0;
    assign process_intf_5.region_idle = region_1_idle;
    assign process_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;
    df_process_intf process_intf_6(clock,reset);
    assign process_intf_6.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_6.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_ready;
    assign process_intf_6.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_done;
    assign process_intf_6.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_continue;
    assign process_intf_6.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.real_start;
    assign process_intf_6.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_query_1_3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.d_query_1_3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_2_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.d_value_1_3_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.d_query_1_3_blk_n;
    assign process_intf_6.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.k_proj_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.q_proj_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.v_proj_1_blk_n;
    assign process_intf_6.cin_stall = 1'b0;
    assign process_intf_6.cout_stall = 1'b0;
    assign process_intf_6.region_idle = region_1_idle;
    assign process_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_6;
    csv_file_dump pstatus_csv_dumper_6;
    df_process_monitor process_monitor_6;
    df_process_intf process_intf_7(clock,reset);
    assign process_intf_7.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.ap_start;
    assign process_intf_7.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.ap_ready;
    assign process_intf_7.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.ap_done;
    assign process_intf_7.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.ap_continue;
    assign process_intf_7.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.ap_start;
    assign process_intf_7.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.q_proj_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.k_proj_0_blk_n;
    assign process_intf_7.pout_stall = 1'b0;
    assign process_intf_7.cin_stall = 1'b0;
    assign process_intf_7.cout_stall = 1'b0;
    assign process_intf_7.region_idle = region_1_idle;
    assign process_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_7;
    csv_file_dump pstatus_csv_dumper_7;
    df_process_monitor process_monitor_7;
    df_process_intf process_intf_8(clock,reset);
    assign process_intf_8.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.ap_start;
    assign process_intf_8.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.ap_ready;
    assign process_intf_8.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.ap_done;
    assign process_intf_8.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.ap_continue;
    assign process_intf_8.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.ap_start;
    assign process_intf_8.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.q_proj_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.k_proj_1_blk_n;
    assign process_intf_8.pout_stall = 1'b0;
    assign process_intf_8.cin_stall = 1'b0;
    assign process_intf_8.cout_stall = 1'b0;
    assign process_intf_8.region_idle = region_1_idle;
    assign process_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_8;
    csv_file_dump pstatus_csv_dumper_8;
    df_process_monitor process_monitor_8;
    df_process_intf process_intf_9(clock,reset);
    assign process_intf_9.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_start;
    assign process_intf_9.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_ready;
    assign process_intf_9.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_done;
    assign process_intf_9.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.ap_continue;
    assign process_intf_9.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.real_start;
    assign process_intf_9.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.v_proj_0_blk_n;
    assign process_intf_9.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.matr_out_0_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.matr_out_0_1_blk_n;
    assign process_intf_9.cin_stall = 1'b0;
    assign process_intf_9.cout_stall = 1'b0;
    assign process_intf_9.region_idle = region_1_idle;
    assign process_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_9;
    csv_file_dump pstatus_csv_dumper_9;
    df_process_monitor process_monitor_9;
    df_process_intf process_intf_10(clock,reset);
    assign process_intf_10.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_10.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_ready;
    assign process_intf_10.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_done;
    assign process_intf_10.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_continue;
    assign process_intf_10.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_10.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.v_proj_1_blk_n;
    assign process_intf_10.pout_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_1_blk_n;
    assign process_intf_10.cin_stall = 1'b0;
    assign process_intf_10.cout_stall = 1'b0;
    assign process_intf_10.region_idle = region_1_idle;
    assign process_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_10;
    csv_file_dump pstatus_csv_dumper_10;
    df_process_monitor process_monitor_10;
    df_process_intf process_intf_11(clock,reset);
    assign process_intf_11.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_11.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_ready;
    assign process_intf_11.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_done;
    assign process_intf_11.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_continue;
    assign process_intf_11.real_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.ap_start;
    assign process_intf_11.pin_stall = 1'b0 | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_0_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_0_1_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_0_blk_n | ~AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.dense_out_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.matr_out_1_1_blk_n;
    assign process_intf_11.pout_stall = 1'b0;
    assign process_intf_11.cin_stall = 1'b0;
    assign process_intf_11.cout_stall = 1'b0;
    assign process_intf_11.region_idle = region_1_idle;
    assign process_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_11;
    csv_file_dump pstatus_csv_dumper_11;
    df_process_monitor process_monitor_11;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_myproject.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_myproject.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_myproject.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_done;
    assign module_intf_2.ap_continue = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.ap_continue;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_2_fu_97.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_2_fu_97.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_2_fu_97.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_1_fu_109.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_1_fu_109.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_1_fu_109.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_s_fu_121.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_s_fu_121.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_s_fu_121.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_73.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_read_stream_array_ap_fixed_16_6_5_3_0_4_s_fu_85.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_2_fu_97.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_2_fu_97.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_2_fu_97.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_1_fu_109.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_1_fu_109.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_1_fu_109.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_s_fu_121.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_s_fu_121.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.lin_projection_ap_fixed_ap_fixed_16_6_5_3_0_config3_U0.grp_dense_latency_ap_fixed_ap_fixed_16_6_5_3_0_config3_1_s_fu_121.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_50.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_50.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_50.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_78.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_78.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_78.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_106.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_106.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_106.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_134.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_134.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_134.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_162.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_162.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_162.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_190.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_190.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_190.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_218.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_218.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_218.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_246.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_246.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_246.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_274.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_274.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_274.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_302.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_302.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_302.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_330.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_330.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_330.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_358.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_358.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_358.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_386.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_386.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_386.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_414.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_414.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_414.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_442.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_442.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_442.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_470.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_470.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_470.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_498.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_498.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_498.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_526.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_526.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_526.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_554.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_554.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_554.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_582.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_582.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_1_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_582.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_50.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_50.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_50.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_78.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_78.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_78.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_106.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_106.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_106.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_134.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_134.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_134.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_162.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_162.ap_ready;
    assign module_intf_37.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_162.ap_done;
    assign module_intf_37.ap_continue = 1'b1;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_190.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_190.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_190.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_218.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_218.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_218.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_246.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_246.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_246.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_274.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_274.ap_ready;
    assign module_intf_41.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_274.ap_done;
    assign module_intf_41.ap_continue = 1'b1;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_302.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_302.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_302.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_330.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_330.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_330.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_358.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_358.ap_ready;
    assign module_intf_44.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_358.ap_done;
    assign module_intf_44.ap_continue = 1'b1;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_386.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_386.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_386.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_414.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_414.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_414.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_442.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_442.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_442.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_470.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_470.ap_ready;
    assign module_intf_48.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_470.ap_done;
    assign module_intf_48.ap_continue = 1'b1;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_498.ap_start;
    assign module_intf_49.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_498.ap_ready;
    assign module_intf_49.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_498.ap_done;
    assign module_intf_49.ap_continue = 1'b1;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_526.ap_start;
    assign module_intf_50.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_526.ap_ready;
    assign module_intf_50.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_526.ap_done;
    assign module_intf_50.ap_continue = 1'b1;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_554.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_554.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_554.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_582.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_582.ap_ready;
    assign module_intf_52.ap_done = AESL_inst_myproject.grp_multiheadattention_ap_fixed_ap_fixed_config3_s_fu_206.matrixmul_transpose_ap_fixed_ap_fixed_config3_U0.grp_softmax_legacy_ap_fixed_ap_fixed_softmax_config3_s_fu_582.ap_done;
    assign module_intf_52.ap_continue = 1'b1;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = 1'b0;
    assign module_intf_53.ap_ready = 1'b0;
    assign module_intf_53.ap_done = 1'b0;
    assign module_intf_53.ap_continue = 1'b0;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;


    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);
    fifo_csv_dumper_35 = new("./depth35.csv");
    cstatus_csv_dumper_35 = new("./chan_status35.csv");
    fifo_monitor_35 = new(fifo_csv_dumper_35,fifo_intf_35,cstatus_csv_dumper_35);
    fifo_csv_dumper_36 = new("./depth36.csv");
    cstatus_csv_dumper_36 = new("./chan_status36.csv");
    fifo_monitor_36 = new(fifo_csv_dumper_36,fifo_intf_36,cstatus_csv_dumper_36);
    fifo_csv_dumper_37 = new("./depth37.csv");
    cstatus_csv_dumper_37 = new("./chan_status37.csv");
    fifo_monitor_37 = new(fifo_csv_dumper_37,fifo_intf_37,cstatus_csv_dumper_37);
    fifo_csv_dumper_38 = new("./depth38.csv");
    cstatus_csv_dumper_38 = new("./chan_status38.csv");
    fifo_monitor_38 = new(fifo_csv_dumper_38,fifo_intf_38,cstatus_csv_dumper_38);
    fifo_csv_dumper_39 = new("./depth39.csv");
    cstatus_csv_dumper_39 = new("./chan_status39.csv");
    fifo_monitor_39 = new(fifo_csv_dumper_39,fifo_intf_39,cstatus_csv_dumper_39);
    fifo_csv_dumper_40 = new("./depth40.csv");
    cstatus_csv_dumper_40 = new("./chan_status40.csv");
    fifo_monitor_40 = new(fifo_csv_dumper_40,fifo_intf_40,cstatus_csv_dumper_40);
    fifo_csv_dumper_41 = new("./depth41.csv");
    cstatus_csv_dumper_41 = new("./chan_status41.csv");
    fifo_monitor_41 = new(fifo_csv_dumper_41,fifo_intf_41,cstatus_csv_dumper_41);
    fifo_csv_dumper_42 = new("./depth42.csv");
    cstatus_csv_dumper_42 = new("./chan_status42.csv");
    fifo_monitor_42 = new(fifo_csv_dumper_42,fifo_intf_42,cstatus_csv_dumper_42);
    fifo_csv_dumper_43 = new("./depth43.csv");
    cstatus_csv_dumper_43 = new("./chan_status43.csv");
    fifo_monitor_43 = new(fifo_csv_dumper_43,fifo_intf_43,cstatus_csv_dumper_43);
    fifo_csv_dumper_44 = new("./depth44.csv");
    cstatus_csv_dumper_44 = new("./chan_status44.csv");
    fifo_monitor_44 = new(fifo_csv_dumper_44,fifo_intf_44,cstatus_csv_dumper_44);
    fifo_csv_dumper_45 = new("./depth45.csv");
    cstatus_csv_dumper_45 = new("./chan_status45.csv");
    fifo_monitor_45 = new(fifo_csv_dumper_45,fifo_intf_45,cstatus_csv_dumper_45);
    fifo_csv_dumper_46 = new("./depth46.csv");
    cstatus_csv_dumper_46 = new("./chan_status46.csv");
    fifo_monitor_46 = new(fifo_csv_dumper_46,fifo_intf_46,cstatus_csv_dumper_46);
    fifo_csv_dumper_47 = new("./depth47.csv");
    cstatus_csv_dumper_47 = new("./chan_status47.csv");
    fifo_monitor_47 = new(fifo_csv_dumper_47,fifo_intf_47,cstatus_csv_dumper_47);
    fifo_csv_dumper_48 = new("./depth48.csv");
    cstatus_csv_dumper_48 = new("./chan_status48.csv");
    fifo_monitor_48 = new(fifo_csv_dumper_48,fifo_intf_48,cstatus_csv_dumper_48);
    fifo_csv_dumper_49 = new("./depth49.csv");
    cstatus_csv_dumper_49 = new("./chan_status49.csv");
    fifo_monitor_49 = new(fifo_csv_dumper_49,fifo_intf_49,cstatus_csv_dumper_49);
    fifo_csv_dumper_50 = new("./depth50.csv");
    cstatus_csv_dumper_50 = new("./chan_status50.csv");
    fifo_monitor_50 = new(fifo_csv_dumper_50,fifo_intf_50,cstatus_csv_dumper_50);
    fifo_csv_dumper_51 = new("./depth51.csv");
    cstatus_csv_dumper_51 = new("./chan_status51.csv");
    fifo_monitor_51 = new(fifo_csv_dumper_51,fifo_intf_51,cstatus_csv_dumper_51);
    fifo_csv_dumper_52 = new("./depth52.csv");
    cstatus_csv_dumper_52 = new("./chan_status52.csv");
    fifo_monitor_52 = new(fifo_csv_dumper_52,fifo_intf_52,cstatus_csv_dumper_52);
    fifo_csv_dumper_53 = new("./depth53.csv");
    cstatus_csv_dumper_53 = new("./chan_status53.csv");
    fifo_monitor_53 = new(fifo_csv_dumper_53,fifo_intf_53,cstatus_csv_dumper_53);
    fifo_csv_dumper_54 = new("./depth54.csv");
    cstatus_csv_dumper_54 = new("./chan_status54.csv");
    fifo_monitor_54 = new(fifo_csv_dumper_54,fifo_intf_54,cstatus_csv_dumper_54);
    fifo_csv_dumper_55 = new("./depth55.csv");
    cstatus_csv_dumper_55 = new("./chan_status55.csv");
    fifo_monitor_55 = new(fifo_csv_dumper_55,fifo_intf_55,cstatus_csv_dumper_55);
    fifo_csv_dumper_56 = new("./depth56.csv");
    cstatus_csv_dumper_56 = new("./chan_status56.csv");
    fifo_monitor_56 = new(fifo_csv_dumper_56,fifo_intf_56,cstatus_csv_dumper_56);
    fifo_csv_dumper_57 = new("./depth57.csv");
    cstatus_csv_dumper_57 = new("./chan_status57.csv");
    fifo_monitor_57 = new(fifo_csv_dumper_57,fifo_intf_57,cstatus_csv_dumper_57);
    fifo_csv_dumper_58 = new("./depth58.csv");
    cstatus_csv_dumper_58 = new("./chan_status58.csv");
    fifo_monitor_58 = new(fifo_csv_dumper_58,fifo_intf_58,cstatus_csv_dumper_58);
    fifo_csv_dumper_59 = new("./depth59.csv");
    cstatus_csv_dumper_59 = new("./chan_status59.csv");
    fifo_monitor_59 = new(fifo_csv_dumper_59,fifo_intf_59,cstatus_csv_dumper_59);
    fifo_csv_dumper_60 = new("./depth60.csv");
    cstatus_csv_dumper_60 = new("./chan_status60.csv");
    fifo_monitor_60 = new(fifo_csv_dumper_60,fifo_intf_60,cstatus_csv_dumper_60);
    fifo_csv_dumper_61 = new("./depth61.csv");
    cstatus_csv_dumper_61 = new("./chan_status61.csv");
    fifo_monitor_61 = new(fifo_csv_dumper_61,fifo_intf_61,cstatus_csv_dumper_61);
    fifo_csv_dumper_62 = new("./depth62.csv");
    cstatus_csv_dumper_62 = new("./chan_status62.csv");
    fifo_monitor_62 = new(fifo_csv_dumper_62,fifo_intf_62,cstatus_csv_dumper_62);
    fifo_csv_dumper_63 = new("./depth63.csv");
    cstatus_csv_dumper_63 = new("./chan_status63.csv");
    fifo_monitor_63 = new(fifo_csv_dumper_63,fifo_intf_63,cstatus_csv_dumper_63);
    fifo_csv_dumper_64 = new("./depth64.csv");
    cstatus_csv_dumper_64 = new("./chan_status64.csv");
    fifo_monitor_64 = new(fifo_csv_dumper_64,fifo_intf_64,cstatus_csv_dumper_64);
    fifo_csv_dumper_65 = new("./depth65.csv");
    cstatus_csv_dumper_65 = new("./chan_status65.csv");
    fifo_monitor_65 = new(fifo_csv_dumper_65,fifo_intf_65,cstatus_csv_dumper_65);
    fifo_csv_dumper_66 = new("./depth66.csv");
    cstatus_csv_dumper_66 = new("./chan_status66.csv");
    fifo_monitor_66 = new(fifo_csv_dumper_66,fifo_intf_66,cstatus_csv_dumper_66);
    fifo_csv_dumper_67 = new("./depth67.csv");
    cstatus_csv_dumper_67 = new("./chan_status67.csv");
    fifo_monitor_67 = new(fifo_csv_dumper_67,fifo_intf_67,cstatus_csv_dumper_67);
    fifo_csv_dumper_68 = new("./depth68.csv");
    cstatus_csv_dumper_68 = new("./chan_status68.csv");
    fifo_monitor_68 = new(fifo_csv_dumper_68,fifo_intf_68,cstatus_csv_dumper_68);
    fifo_csv_dumper_69 = new("./depth69.csv");
    cstatus_csv_dumper_69 = new("./chan_status69.csv");
    fifo_monitor_69 = new(fifo_csv_dumper_69,fifo_intf_69,cstatus_csv_dumper_69);
    fifo_csv_dumper_70 = new("./depth70.csv");
    cstatus_csv_dumper_70 = new("./chan_status70.csv");
    fifo_monitor_70 = new(fifo_csv_dumper_70,fifo_intf_70,cstatus_csv_dumper_70);
    fifo_csv_dumper_71 = new("./depth71.csv");
    cstatus_csv_dumper_71 = new("./chan_status71.csv");
    fifo_monitor_71 = new(fifo_csv_dumper_71,fifo_intf_71,cstatus_csv_dumper_71);
    fifo_csv_dumper_72 = new("./depth72.csv");
    cstatus_csv_dumper_72 = new("./chan_status72.csv");
    fifo_monitor_72 = new(fifo_csv_dumper_72,fifo_intf_72,cstatus_csv_dumper_72);
    fifo_csv_dumper_73 = new("./depth73.csv");
    cstatus_csv_dumper_73 = new("./chan_status73.csv");
    fifo_monitor_73 = new(fifo_csv_dumper_73,fifo_intf_73,cstatus_csv_dumper_73);
    fifo_csv_dumper_74 = new("./depth74.csv");
    cstatus_csv_dumper_74 = new("./chan_status74.csv");
    fifo_monitor_74 = new(fifo_csv_dumper_74,fifo_intf_74,cstatus_csv_dumper_74);
    fifo_csv_dumper_75 = new("./depth75.csv");
    cstatus_csv_dumper_75 = new("./chan_status75.csv");
    fifo_monitor_75 = new(fifo_csv_dumper_75,fifo_intf_75,cstatus_csv_dumper_75);
    fifo_csv_dumper_76 = new("./depth76.csv");
    cstatus_csv_dumper_76 = new("./chan_status76.csv");
    fifo_monitor_76 = new(fifo_csv_dumper_76,fifo_intf_76,cstatus_csv_dumper_76);
    fifo_csv_dumper_77 = new("./depth77.csv");
    cstatus_csv_dumper_77 = new("./chan_status77.csv");
    fifo_monitor_77 = new(fifo_csv_dumper_77,fifo_intf_77,cstatus_csv_dumper_77);
    fifo_csv_dumper_78 = new("./depth78.csv");
    cstatus_csv_dumper_78 = new("./chan_status78.csv");
    fifo_monitor_78 = new(fifo_csv_dumper_78,fifo_intf_78,cstatus_csv_dumper_78);
    fifo_csv_dumper_79 = new("./depth79.csv");
    cstatus_csv_dumper_79 = new("./chan_status79.csv");
    fifo_monitor_79 = new(fifo_csv_dumper_79,fifo_intf_79,cstatus_csv_dumper_79);
    fifo_csv_dumper_80 = new("./depth80.csv");
    cstatus_csv_dumper_80 = new("./chan_status80.csv");
    fifo_monitor_80 = new(fifo_csv_dumper_80,fifo_intf_80,cstatus_csv_dumper_80);
    fifo_csv_dumper_81 = new("./depth81.csv");
    cstatus_csv_dumper_81 = new("./chan_status81.csv");
    fifo_monitor_81 = new(fifo_csv_dumper_81,fifo_intf_81,cstatus_csv_dumper_81);
    fifo_csv_dumper_82 = new("./depth82.csv");
    cstatus_csv_dumper_82 = new("./chan_status82.csv");
    fifo_monitor_82 = new(fifo_csv_dumper_82,fifo_intf_82,cstatus_csv_dumper_82);
    fifo_csv_dumper_83 = new("./depth83.csv");
    cstatus_csv_dumper_83 = new("./chan_status83.csv");
    fifo_monitor_83 = new(fifo_csv_dumper_83,fifo_intf_83,cstatus_csv_dumper_83);
    fifo_csv_dumper_84 = new("./depth84.csv");
    cstatus_csv_dumper_84 = new("./chan_status84.csv");
    fifo_monitor_84 = new(fifo_csv_dumper_84,fifo_intf_84,cstatus_csv_dumper_84);
    fifo_csv_dumper_85 = new("./depth85.csv");
    cstatus_csv_dumper_85 = new("./chan_status85.csv");
    fifo_monitor_85 = new(fifo_csv_dumper_85,fifo_intf_85,cstatus_csv_dumper_85);
    fifo_csv_dumper_86 = new("./depth86.csv");
    cstatus_csv_dumper_86 = new("./chan_status86.csv");
    fifo_monitor_86 = new(fifo_csv_dumper_86,fifo_intf_86,cstatus_csv_dumper_86);
    fifo_csv_dumper_87 = new("./depth87.csv");
    cstatus_csv_dumper_87 = new("./chan_status87.csv");
    fifo_monitor_87 = new(fifo_csv_dumper_87,fifo_intf_87,cstatus_csv_dumper_87);
    fifo_csv_dumper_88 = new("./depth88.csv");
    cstatus_csv_dumper_88 = new("./chan_status88.csv");
    fifo_monitor_88 = new(fifo_csv_dumper_88,fifo_intf_88,cstatus_csv_dumper_88);
    fifo_csv_dumper_89 = new("./depth89.csv");
    cstatus_csv_dumper_89 = new("./chan_status89.csv");
    fifo_monitor_89 = new(fifo_csv_dumper_89,fifo_intf_89,cstatus_csv_dumper_89);
    fifo_csv_dumper_90 = new("./depth90.csv");
    cstatus_csv_dumper_90 = new("./chan_status90.csv");
    fifo_monitor_90 = new(fifo_csv_dumper_90,fifo_intf_90,cstatus_csv_dumper_90);
    fifo_csv_dumper_91 = new("./depth91.csv");
    cstatus_csv_dumper_91 = new("./chan_status91.csv");
    fifo_monitor_91 = new(fifo_csv_dumper_91,fifo_intf_91,cstatus_csv_dumper_91);
    fifo_csv_dumper_92 = new("./depth92.csv");
    cstatus_csv_dumper_92 = new("./chan_status92.csv");
    fifo_monitor_92 = new(fifo_csv_dumper_92,fifo_intf_92,cstatus_csv_dumper_92);
    fifo_csv_dumper_93 = new("./depth93.csv");
    cstatus_csv_dumper_93 = new("./chan_status93.csv");
    fifo_monitor_93 = new(fifo_csv_dumper_93,fifo_intf_93,cstatus_csv_dumper_93);
    fifo_csv_dumper_94 = new("./depth94.csv");
    cstatus_csv_dumper_94 = new("./chan_status94.csv");
    fifo_monitor_94 = new(fifo_csv_dumper_94,fifo_intf_94,cstatus_csv_dumper_94);
    fifo_csv_dumper_95 = new("./depth95.csv");
    cstatus_csv_dumper_95 = new("./chan_status95.csv");
    fifo_monitor_95 = new(fifo_csv_dumper_95,fifo_intf_95,cstatus_csv_dumper_95);
    fifo_csv_dumper_96 = new("./depth96.csv");
    cstatus_csv_dumper_96 = new("./chan_status96.csv");
    fifo_monitor_96 = new(fifo_csv_dumper_96,fifo_intf_96,cstatus_csv_dumper_96);
    fifo_csv_dumper_97 = new("./depth97.csv");
    cstatus_csv_dumper_97 = new("./chan_status97.csv");
    fifo_monitor_97 = new(fifo_csv_dumper_97,fifo_intf_97,cstatus_csv_dumper_97);
    fifo_csv_dumper_98 = new("./depth98.csv");
    cstatus_csv_dumper_98 = new("./chan_status98.csv");
    fifo_monitor_98 = new(fifo_csv_dumper_98,fifo_intf_98,cstatus_csv_dumper_98);
    fifo_csv_dumper_99 = new("./depth99.csv");
    cstatus_csv_dumper_99 = new("./chan_status99.csv");
    fifo_monitor_99 = new(fifo_csv_dumper_99,fifo_intf_99,cstatus_csv_dumper_99);
    fifo_csv_dumper_100 = new("./depth100.csv");
    cstatus_csv_dumper_100 = new("./chan_status100.csv");
    fifo_monitor_100 = new(fifo_csv_dumper_100,fifo_intf_100,cstatus_csv_dumper_100);
    fifo_csv_dumper_101 = new("./depth101.csv");
    cstatus_csv_dumper_101 = new("./chan_status101.csv");
    fifo_monitor_101 = new(fifo_csv_dumper_101,fifo_intf_101,cstatus_csv_dumper_101);
    fifo_csv_dumper_102 = new("./depth102.csv");
    cstatus_csv_dumper_102 = new("./chan_status102.csv");
    fifo_monitor_102 = new(fifo_csv_dumper_102,fifo_intf_102,cstatus_csv_dumper_102);
    fifo_csv_dumper_103 = new("./depth103.csv");
    cstatus_csv_dumper_103 = new("./chan_status103.csv");
    fifo_monitor_103 = new(fifo_csv_dumper_103,fifo_intf_103,cstatus_csv_dumper_103);
    fifo_csv_dumper_104 = new("./depth104.csv");
    cstatus_csv_dumper_104 = new("./chan_status104.csv");
    fifo_monitor_104 = new(fifo_csv_dumper_104,fifo_intf_104,cstatus_csv_dumper_104);
    fifo_csv_dumper_105 = new("./depth105.csv");
    cstatus_csv_dumper_105 = new("./chan_status105.csv");
    fifo_monitor_105 = new(fifo_csv_dumper_105,fifo_intf_105,cstatus_csv_dumper_105);
    fifo_csv_dumper_106 = new("./depth106.csv");
    cstatus_csv_dumper_106 = new("./chan_status106.csv");
    fifo_monitor_106 = new(fifo_csv_dumper_106,fifo_intf_106,cstatus_csv_dumper_106);
    fifo_csv_dumper_107 = new("./depth107.csv");
    cstatus_csv_dumper_107 = new("./chan_status107.csv");
    fifo_monitor_107 = new(fifo_csv_dumper_107,fifo_intf_107,cstatus_csv_dumper_107);
    fifo_csv_dumper_108 = new("./depth108.csv");
    cstatus_csv_dumper_108 = new("./chan_status108.csv");
    fifo_monitor_108 = new(fifo_csv_dumper_108,fifo_intf_108,cstatus_csv_dumper_108);
    fifo_csv_dumper_109 = new("./depth109.csv");
    cstatus_csv_dumper_109 = new("./chan_status109.csv");
    fifo_monitor_109 = new(fifo_csv_dumper_109,fifo_intf_109,cstatus_csv_dumper_109);
    fifo_csv_dumper_110 = new("./depth110.csv");
    cstatus_csv_dumper_110 = new("./chan_status110.csv");
    fifo_monitor_110 = new(fifo_csv_dumper_110,fifo_intf_110,cstatus_csv_dumper_110);
    fifo_csv_dumper_111 = new("./depth111.csv");
    cstatus_csv_dumper_111 = new("./chan_status111.csv");
    fifo_monitor_111 = new(fifo_csv_dumper_111,fifo_intf_111,cstatus_csv_dumper_111);
    fifo_csv_dumper_112 = new("./depth112.csv");
    cstatus_csv_dumper_112 = new("./chan_status112.csv");
    fifo_monitor_112 = new(fifo_csv_dumper_112,fifo_intf_112,cstatus_csv_dumper_112);
    fifo_csv_dumper_113 = new("./depth113.csv");
    cstatus_csv_dumper_113 = new("./chan_status113.csv");
    fifo_monitor_113 = new(fifo_csv_dumper_113,fifo_intf_113,cstatus_csv_dumper_113);
    fifo_csv_dumper_114 = new("./depth114.csv");
    cstatus_csv_dumper_114 = new("./chan_status114.csv");
    fifo_monitor_114 = new(fifo_csv_dumper_114,fifo_intf_114,cstatus_csv_dumper_114);
    fifo_csv_dumper_115 = new("./depth115.csv");
    cstatus_csv_dumper_115 = new("./chan_status115.csv");
    fifo_monitor_115 = new(fifo_csv_dumper_115,fifo_intf_115,cstatus_csv_dumper_115);
    fifo_csv_dumper_116 = new("./depth116.csv");
    cstatus_csv_dumper_116 = new("./chan_status116.csv");
    fifo_monitor_116 = new(fifo_csv_dumper_116,fifo_intf_116,cstatus_csv_dumper_116);
    fifo_csv_dumper_117 = new("./depth117.csv");
    cstatus_csv_dumper_117 = new("./chan_status117.csv");
    fifo_monitor_117 = new(fifo_csv_dumper_117,fifo_intf_117,cstatus_csv_dumper_117);
    fifo_csv_dumper_118 = new("./depth118.csv");
    cstatus_csv_dumper_118 = new("./chan_status118.csv");
    fifo_monitor_118 = new(fifo_csv_dumper_118,fifo_intf_118,cstatus_csv_dumper_118);
    fifo_csv_dumper_119 = new("./depth119.csv");
    cstatus_csv_dumper_119 = new("./chan_status119.csv");
    fifo_monitor_119 = new(fifo_csv_dumper_119,fifo_intf_119,cstatus_csv_dumper_119);
    fifo_csv_dumper_120 = new("./depth120.csv");
    cstatus_csv_dumper_120 = new("./chan_status120.csv");
    fifo_monitor_120 = new(fifo_csv_dumper_120,fifo_intf_120,cstatus_csv_dumper_120);
    fifo_csv_dumper_121 = new("./depth121.csv");
    cstatus_csv_dumper_121 = new("./chan_status121.csv");
    fifo_monitor_121 = new(fifo_csv_dumper_121,fifo_intf_121,cstatus_csv_dumper_121);
    fifo_csv_dumper_122 = new("./depth122.csv");
    cstatus_csv_dumper_122 = new("./chan_status122.csv");
    fifo_monitor_122 = new(fifo_csv_dumper_122,fifo_intf_122,cstatus_csv_dumper_122);
    fifo_csv_dumper_123 = new("./depth123.csv");
    cstatus_csv_dumper_123 = new("./chan_status123.csv");
    fifo_monitor_123 = new(fifo_csv_dumper_123,fifo_intf_123,cstatus_csv_dumper_123);
    fifo_csv_dumper_124 = new("./depth124.csv");
    cstatus_csv_dumper_124 = new("./chan_status124.csv");
    fifo_monitor_124 = new(fifo_csv_dumper_124,fifo_intf_124,cstatus_csv_dumper_124);
    fifo_csv_dumper_125 = new("./depth125.csv");
    cstatus_csv_dumper_125 = new("./chan_status125.csv");
    fifo_monitor_125 = new(fifo_csv_dumper_125,fifo_intf_125,cstatus_csv_dumper_125);
    fifo_csv_dumper_126 = new("./depth126.csv");
    cstatus_csv_dumper_126 = new("./chan_status126.csv");
    fifo_monitor_126 = new(fifo_csv_dumper_126,fifo_intf_126,cstatus_csv_dumper_126);
    fifo_csv_dumper_127 = new("./depth127.csv");
    cstatus_csv_dumper_127 = new("./chan_status127.csv");
    fifo_monitor_127 = new(fifo_csv_dumper_127,fifo_intf_127,cstatus_csv_dumper_127);
    fifo_csv_dumper_128 = new("./depth128.csv");
    cstatus_csv_dumper_128 = new("./chan_status128.csv");
    fifo_monitor_128 = new(fifo_csv_dumper_128,fifo_intf_128,cstatus_csv_dumper_128);
    fifo_csv_dumper_129 = new("./depth129.csv");
    cstatus_csv_dumper_129 = new("./chan_status129.csv");
    fifo_monitor_129 = new(fifo_csv_dumper_129,fifo_intf_129,cstatus_csv_dumper_129);
    fifo_csv_dumper_130 = new("./depth130.csv");
    cstatus_csv_dumper_130 = new("./chan_status130.csv");
    fifo_monitor_130 = new(fifo_csv_dumper_130,fifo_intf_130,cstatus_csv_dumper_130);
    fifo_csv_dumper_131 = new("./depth131.csv");
    cstatus_csv_dumper_131 = new("./chan_status131.csv");
    fifo_monitor_131 = new(fifo_csv_dumper_131,fifo_intf_131,cstatus_csv_dumper_131);
    fifo_csv_dumper_132 = new("./depth132.csv");
    cstatus_csv_dumper_132 = new("./chan_status132.csv");
    fifo_monitor_132 = new(fifo_csv_dumper_132,fifo_intf_132,cstatus_csv_dumper_132);
    fifo_csv_dumper_133 = new("./depth133.csv");
    cstatus_csv_dumper_133 = new("./chan_status133.csv");
    fifo_monitor_133 = new(fifo_csv_dumper_133,fifo_intf_133,cstatus_csv_dumper_133);
    fifo_csv_dumper_134 = new("./depth134.csv");
    cstatus_csv_dumper_134 = new("./chan_status134.csv");
    fifo_monitor_134 = new(fifo_csv_dumper_134,fifo_intf_134,cstatus_csv_dumper_134);
    fifo_csv_dumper_135 = new("./depth135.csv");
    cstatus_csv_dumper_135 = new("./chan_status135.csv");
    fifo_monitor_135 = new(fifo_csv_dumper_135,fifo_intf_135,cstatus_csv_dumper_135);
    fifo_csv_dumper_136 = new("./depth136.csv");
    cstatus_csv_dumper_136 = new("./chan_status136.csv");
    fifo_monitor_136 = new(fifo_csv_dumper_136,fifo_intf_136,cstatus_csv_dumper_136);
    fifo_csv_dumper_137 = new("./depth137.csv");
    cstatus_csv_dumper_137 = new("./chan_status137.csv");
    fifo_monitor_137 = new(fifo_csv_dumper_137,fifo_intf_137,cstatus_csv_dumper_137);
    fifo_csv_dumper_138 = new("./depth138.csv");
    cstatus_csv_dumper_138 = new("./chan_status138.csv");
    fifo_monitor_138 = new(fifo_csv_dumper_138,fifo_intf_138,cstatus_csv_dumper_138);
    fifo_csv_dumper_139 = new("./depth139.csv");
    cstatus_csv_dumper_139 = new("./chan_status139.csv");
    fifo_monitor_139 = new(fifo_csv_dumper_139,fifo_intf_139,cstatus_csv_dumper_139);
    fifo_csv_dumper_140 = new("./depth140.csv");
    cstatus_csv_dumper_140 = new("./chan_status140.csv");
    fifo_monitor_140 = new(fifo_csv_dumper_140,fifo_intf_140,cstatus_csv_dumper_140);
    fifo_csv_dumper_141 = new("./depth141.csv");
    cstatus_csv_dumper_141 = new("./chan_status141.csv");
    fifo_monitor_141 = new(fifo_csv_dumper_141,fifo_intf_141,cstatus_csv_dumper_141);
    fifo_csv_dumper_142 = new("./depth142.csv");
    cstatus_csv_dumper_142 = new("./chan_status142.csv");
    fifo_monitor_142 = new(fifo_csv_dumper_142,fifo_intf_142,cstatus_csv_dumper_142);
    fifo_csv_dumper_143 = new("./depth143.csv");
    cstatus_csv_dumper_143 = new("./chan_status143.csv");
    fifo_monitor_143 = new(fifo_csv_dumper_143,fifo_intf_143,cstatus_csv_dumper_143);
    fifo_csv_dumper_144 = new("./depth144.csv");
    cstatus_csv_dumper_144 = new("./chan_status144.csv");
    fifo_monitor_144 = new(fifo_csv_dumper_144,fifo_intf_144,cstatus_csv_dumper_144);
    fifo_csv_dumper_145 = new("./depth145.csv");
    cstatus_csv_dumper_145 = new("./chan_status145.csv");
    fifo_monitor_145 = new(fifo_csv_dumper_145,fifo_intf_145,cstatus_csv_dumper_145);
    fifo_csv_dumper_146 = new("./depth146.csv");
    cstatus_csv_dumper_146 = new("./chan_status146.csv");
    fifo_monitor_146 = new(fifo_csv_dumper_146,fifo_intf_146,cstatus_csv_dumper_146);
    fifo_csv_dumper_147 = new("./depth147.csv");
    cstatus_csv_dumper_147 = new("./chan_status147.csv");
    fifo_monitor_147 = new(fifo_csv_dumper_147,fifo_intf_147,cstatus_csv_dumper_147);
    fifo_csv_dumper_148 = new("./depth148.csv");
    cstatus_csv_dumper_148 = new("./chan_status148.csv");
    fifo_monitor_148 = new(fifo_csv_dumper_148,fifo_intf_148,cstatus_csv_dumper_148);
    fifo_csv_dumper_149 = new("./depth149.csv");
    cstatus_csv_dumper_149 = new("./chan_status149.csv");
    fifo_monitor_149 = new(fifo_csv_dumper_149,fifo_intf_149,cstatus_csv_dumper_149);
    fifo_csv_dumper_150 = new("./depth150.csv");
    cstatus_csv_dumper_150 = new("./chan_status150.csv");
    fifo_monitor_150 = new(fifo_csv_dumper_150,fifo_intf_150,cstatus_csv_dumper_150);
    fifo_csv_dumper_151 = new("./depth151.csv");
    cstatus_csv_dumper_151 = new("./chan_status151.csv");
    fifo_monitor_151 = new(fifo_csv_dumper_151,fifo_intf_151,cstatus_csv_dumper_151);
    fifo_csv_dumper_152 = new("./depth152.csv");
    cstatus_csv_dumper_152 = new("./chan_status152.csv");
    fifo_monitor_152 = new(fifo_csv_dumper_152,fifo_intf_152,cstatus_csv_dumper_152);
    fifo_csv_dumper_153 = new("./depth153.csv");
    cstatus_csv_dumper_153 = new("./chan_status153.csv");
    fifo_monitor_153 = new(fifo_csv_dumper_153,fifo_intf_153,cstatus_csv_dumper_153);
    fifo_csv_dumper_154 = new("./depth154.csv");
    cstatus_csv_dumper_154 = new("./chan_status154.csv");
    fifo_monitor_154 = new(fifo_csv_dumper_154,fifo_intf_154,cstatus_csv_dumper_154);
    fifo_csv_dumper_155 = new("./depth155.csv");
    cstatus_csv_dumper_155 = new("./chan_status155.csv");
    fifo_monitor_155 = new(fifo_csv_dumper_155,fifo_intf_155,cstatus_csv_dumper_155);
    fifo_csv_dumper_156 = new("./depth156.csv");
    cstatus_csv_dumper_156 = new("./chan_status156.csv");
    fifo_monitor_156 = new(fifo_csv_dumper_156,fifo_intf_156,cstatus_csv_dumper_156);
    fifo_csv_dumper_157 = new("./depth157.csv");
    cstatus_csv_dumper_157 = new("./chan_status157.csv");
    fifo_monitor_157 = new(fifo_csv_dumper_157,fifo_intf_157,cstatus_csv_dumper_157);
    fifo_csv_dumper_158 = new("./depth158.csv");
    cstatus_csv_dumper_158 = new("./chan_status158.csv");
    fifo_monitor_158 = new(fifo_csv_dumper_158,fifo_intf_158,cstatus_csv_dumper_158);
    fifo_csv_dumper_159 = new("./depth159.csv");
    cstatus_csv_dumper_159 = new("./chan_status159.csv");
    fifo_monitor_159 = new(fifo_csv_dumper_159,fifo_intf_159,cstatus_csv_dumper_159);
    fifo_csv_dumper_160 = new("./depth160.csv");
    cstatus_csv_dumper_160 = new("./chan_status160.csv");
    fifo_monitor_160 = new(fifo_csv_dumper_160,fifo_intf_160,cstatus_csv_dumper_160);
    fifo_csv_dumper_161 = new("./depth161.csv");
    cstatus_csv_dumper_161 = new("./chan_status161.csv");
    fifo_monitor_161 = new(fifo_csv_dumper_161,fifo_intf_161,cstatus_csv_dumper_161);
    fifo_csv_dumper_162 = new("./depth162.csv");
    cstatus_csv_dumper_162 = new("./chan_status162.csv");
    fifo_monitor_162 = new(fifo_csv_dumper_162,fifo_intf_162,cstatus_csv_dumper_162);
    fifo_csv_dumper_163 = new("./depth163.csv");
    cstatus_csv_dumper_163 = new("./chan_status163.csv");
    fifo_monitor_163 = new(fifo_csv_dumper_163,fifo_intf_163,cstatus_csv_dumper_163);
    fifo_csv_dumper_164 = new("./depth164.csv");
    cstatus_csv_dumper_164 = new("./chan_status164.csv");
    fifo_monitor_164 = new(fifo_csv_dumper_164,fifo_intf_164,cstatus_csv_dumper_164);
    fifo_csv_dumper_165 = new("./depth165.csv");
    cstatus_csv_dumper_165 = new("./chan_status165.csv");
    fifo_monitor_165 = new(fifo_csv_dumper_165,fifo_intf_165,cstatus_csv_dumper_165);
    fifo_csv_dumper_166 = new("./depth166.csv");
    cstatus_csv_dumper_166 = new("./chan_status166.csv");
    fifo_monitor_166 = new(fifo_csv_dumper_166,fifo_intf_166,cstatus_csv_dumper_166);
    fifo_csv_dumper_167 = new("./depth167.csv");
    cstatus_csv_dumper_167 = new("./chan_status167.csv");
    fifo_monitor_167 = new(fifo_csv_dumper_167,fifo_intf_167,cstatus_csv_dumper_167);
    fifo_csv_dumper_168 = new("./depth168.csv");
    cstatus_csv_dumper_168 = new("./chan_status168.csv");
    fifo_monitor_168 = new(fifo_csv_dumper_168,fifo_intf_168,cstatus_csv_dumper_168);
    fifo_csv_dumper_169 = new("./depth169.csv");
    cstatus_csv_dumper_169 = new("./chan_status169.csv");
    fifo_monitor_169 = new(fifo_csv_dumper_169,fifo_intf_169,cstatus_csv_dumper_169);
    fifo_csv_dumper_170 = new("./depth170.csv");
    cstatus_csv_dumper_170 = new("./chan_status170.csv");
    fifo_monitor_170 = new(fifo_csv_dumper_170,fifo_intf_170,cstatus_csv_dumper_170);
    fifo_csv_dumper_171 = new("./depth171.csv");
    cstatus_csv_dumper_171 = new("./chan_status171.csv");
    fifo_monitor_171 = new(fifo_csv_dumper_171,fifo_intf_171,cstatus_csv_dumper_171);
    fifo_csv_dumper_172 = new("./depth172.csv");
    cstatus_csv_dumper_172 = new("./chan_status172.csv");
    fifo_monitor_172 = new(fifo_csv_dumper_172,fifo_intf_172,cstatus_csv_dumper_172);
    fifo_csv_dumper_173 = new("./depth173.csv");
    cstatus_csv_dumper_173 = new("./chan_status173.csv");
    fifo_monitor_173 = new(fifo_csv_dumper_173,fifo_intf_173,cstatus_csv_dumper_173);
    fifo_csv_dumper_174 = new("./depth174.csv");
    cstatus_csv_dumper_174 = new("./chan_status174.csv");
    fifo_monitor_174 = new(fifo_csv_dumper_174,fifo_intf_174,cstatus_csv_dumper_174);
    fifo_csv_dumper_175 = new("./depth175.csv");
    cstatus_csv_dumper_175 = new("./chan_status175.csv");
    fifo_monitor_175 = new(fifo_csv_dumper_175,fifo_intf_175,cstatus_csv_dumper_175);
    fifo_csv_dumper_176 = new("./depth176.csv");
    cstatus_csv_dumper_176 = new("./chan_status176.csv");
    fifo_monitor_176 = new(fifo_csv_dumper_176,fifo_intf_176,cstatus_csv_dumper_176);
    fifo_csv_dumper_177 = new("./depth177.csv");
    cstatus_csv_dumper_177 = new("./chan_status177.csv");
    fifo_monitor_177 = new(fifo_csv_dumper_177,fifo_intf_177,cstatus_csv_dumper_177);
    fifo_csv_dumper_178 = new("./depth178.csv");
    cstatus_csv_dumper_178 = new("./chan_status178.csv");
    fifo_monitor_178 = new(fifo_csv_dumper_178,fifo_intf_178,cstatus_csv_dumper_178);
    fifo_csv_dumper_179 = new("./depth179.csv");
    cstatus_csv_dumper_179 = new("./chan_status179.csv");
    fifo_monitor_179 = new(fifo_csv_dumper_179,fifo_intf_179,cstatus_csv_dumper_179);
    fifo_csv_dumper_180 = new("./depth180.csv");
    cstatus_csv_dumper_180 = new("./chan_status180.csv");
    fifo_monitor_180 = new(fifo_csv_dumper_180,fifo_intf_180,cstatus_csv_dumper_180);
    fifo_csv_dumper_181 = new("./depth181.csv");
    cstatus_csv_dumper_181 = new("./chan_status181.csv");
    fifo_monitor_181 = new(fifo_csv_dumper_181,fifo_intf_181,cstatus_csv_dumper_181);
    fifo_csv_dumper_182 = new("./depth182.csv");
    cstatus_csv_dumper_182 = new("./chan_status182.csv");
    fifo_monitor_182 = new(fifo_csv_dumper_182,fifo_intf_182,cstatus_csv_dumper_182);
    fifo_csv_dumper_183 = new("./depth183.csv");
    cstatus_csv_dumper_183 = new("./chan_status183.csv");
    fifo_monitor_183 = new(fifo_csv_dumper_183,fifo_intf_183,cstatus_csv_dumper_183);
    fifo_csv_dumper_184 = new("./depth184.csv");
    cstatus_csv_dumper_184 = new("./chan_status184.csv");
    fifo_monitor_184 = new(fifo_csv_dumper_184,fifo_intf_184,cstatus_csv_dumper_184);
    fifo_csv_dumper_185 = new("./depth185.csv");
    cstatus_csv_dumper_185 = new("./chan_status185.csv");
    fifo_monitor_185 = new(fifo_csv_dumper_185,fifo_intf_185,cstatus_csv_dumper_185);
    fifo_csv_dumper_186 = new("./depth186.csv");
    cstatus_csv_dumper_186 = new("./chan_status186.csv");
    fifo_monitor_186 = new(fifo_csv_dumper_186,fifo_intf_186,cstatus_csv_dumper_186);
    fifo_csv_dumper_187 = new("./depth187.csv");
    cstatus_csv_dumper_187 = new("./chan_status187.csv");
    fifo_monitor_187 = new(fifo_csv_dumper_187,fifo_intf_187,cstatus_csv_dumper_187);
    fifo_csv_dumper_188 = new("./depth188.csv");
    cstatus_csv_dumper_188 = new("./chan_status188.csv");
    fifo_monitor_188 = new(fifo_csv_dumper_188,fifo_intf_188,cstatus_csv_dumper_188);
    fifo_csv_dumper_189 = new("./depth189.csv");
    cstatus_csv_dumper_189 = new("./chan_status189.csv");
    fifo_monitor_189 = new(fifo_csv_dumper_189,fifo_intf_189,cstatus_csv_dumper_189);
    fifo_csv_dumper_190 = new("./depth190.csv");
    cstatus_csv_dumper_190 = new("./chan_status190.csv");
    fifo_monitor_190 = new(fifo_csv_dumper_190,fifo_intf_190,cstatus_csv_dumper_190);
    fifo_csv_dumper_191 = new("./depth191.csv");
    cstatus_csv_dumper_191 = new("./chan_status191.csv");
    fifo_monitor_191 = new(fifo_csv_dumper_191,fifo_intf_191,cstatus_csv_dumper_191);
    fifo_csv_dumper_192 = new("./depth192.csv");
    cstatus_csv_dumper_192 = new("./chan_status192.csv");
    fifo_monitor_192 = new(fifo_csv_dumper_192,fifo_intf_192,cstatus_csv_dumper_192);
    fifo_csv_dumper_193 = new("./depth193.csv");
    cstatus_csv_dumper_193 = new("./chan_status193.csv");
    fifo_monitor_193 = new(fifo_csv_dumper_193,fifo_intf_193,cstatus_csv_dumper_193);
    fifo_csv_dumper_194 = new("./depth194.csv");
    cstatus_csv_dumper_194 = new("./chan_status194.csv");
    fifo_monitor_194 = new(fifo_csv_dumper_194,fifo_intf_194,cstatus_csv_dumper_194);
    fifo_csv_dumper_195 = new("./depth195.csv");
    cstatus_csv_dumper_195 = new("./chan_status195.csv");
    fifo_monitor_195 = new(fifo_csv_dumper_195,fifo_intf_195,cstatus_csv_dumper_195);
    fifo_csv_dumper_196 = new("./depth196.csv");
    cstatus_csv_dumper_196 = new("./chan_status196.csv");
    fifo_monitor_196 = new(fifo_csv_dumper_196,fifo_intf_196,cstatus_csv_dumper_196);
    fifo_csv_dumper_197 = new("./depth197.csv");
    cstatus_csv_dumper_197 = new("./chan_status197.csv");
    fifo_monitor_197 = new(fifo_csv_dumper_197,fifo_intf_197,cstatus_csv_dumper_197);
    fifo_csv_dumper_198 = new("./depth198.csv");
    cstatus_csv_dumper_198 = new("./chan_status198.csv");
    fifo_monitor_198 = new(fifo_csv_dumper_198,fifo_intf_198,cstatus_csv_dumper_198);
    fifo_csv_dumper_199 = new("./depth199.csv");
    cstatus_csv_dumper_199 = new("./chan_status199.csv");
    fifo_monitor_199 = new(fifo_csv_dumper_199,fifo_intf_199,cstatus_csv_dumper_199);
    fifo_csv_dumper_200 = new("./depth200.csv");
    cstatus_csv_dumper_200 = new("./chan_status200.csv");
    fifo_monitor_200 = new(fifo_csv_dumper_200,fifo_intf_200,cstatus_csv_dumper_200);
    fifo_csv_dumper_201 = new("./depth201.csv");
    cstatus_csv_dumper_201 = new("./chan_status201.csv");
    fifo_monitor_201 = new(fifo_csv_dumper_201,fifo_intf_201,cstatus_csv_dumper_201);
    fifo_csv_dumper_202 = new("./depth202.csv");
    cstatus_csv_dumper_202 = new("./chan_status202.csv");
    fifo_monitor_202 = new(fifo_csv_dumper_202,fifo_intf_202,cstatus_csv_dumper_202);
    fifo_csv_dumper_203 = new("./depth203.csv");
    cstatus_csv_dumper_203 = new("./chan_status203.csv");
    fifo_monitor_203 = new(fifo_csv_dumper_203,fifo_intf_203,cstatus_csv_dumper_203);
    fifo_csv_dumper_204 = new("./depth204.csv");
    cstatus_csv_dumper_204 = new("./chan_status204.csv");
    fifo_monitor_204 = new(fifo_csv_dumper_204,fifo_intf_204,cstatus_csv_dumper_204);
    fifo_csv_dumper_205 = new("./depth205.csv");
    cstatus_csv_dumper_205 = new("./chan_status205.csv");
    fifo_monitor_205 = new(fifo_csv_dumper_205,fifo_intf_205,cstatus_csv_dumper_205);
    fifo_csv_dumper_206 = new("./depth206.csv");
    cstatus_csv_dumper_206 = new("./chan_status206.csv");
    fifo_monitor_206 = new(fifo_csv_dumper_206,fifo_intf_206,cstatus_csv_dumper_206);
    fifo_csv_dumper_207 = new("./depth207.csv");
    cstatus_csv_dumper_207 = new("./chan_status207.csv");
    fifo_monitor_207 = new(fifo_csv_dumper_207,fifo_intf_207,cstatus_csv_dumper_207);
    fifo_csv_dumper_208 = new("./depth208.csv");
    cstatus_csv_dumper_208 = new("./chan_status208.csv");
    fifo_monitor_208 = new(fifo_csv_dumper_208,fifo_intf_208,cstatus_csv_dumper_208);
    fifo_csv_dumper_209 = new("./depth209.csv");
    cstatus_csv_dumper_209 = new("./chan_status209.csv");
    fifo_monitor_209 = new(fifo_csv_dumper_209,fifo_intf_209,cstatus_csv_dumper_209);
    fifo_csv_dumper_210 = new("./depth210.csv");
    cstatus_csv_dumper_210 = new("./chan_status210.csv");
    fifo_monitor_210 = new(fifo_csv_dumper_210,fifo_intf_210,cstatus_csv_dumper_210);
    fifo_csv_dumper_211 = new("./depth211.csv");
    cstatus_csv_dumper_211 = new("./chan_status211.csv");
    fifo_monitor_211 = new(fifo_csv_dumper_211,fifo_intf_211,cstatus_csv_dumper_211);
    fifo_csv_dumper_212 = new("./depth212.csv");
    cstatus_csv_dumper_212 = new("./chan_status212.csv");
    fifo_monitor_212 = new(fifo_csv_dumper_212,fifo_intf_212,cstatus_csv_dumper_212);
    fifo_csv_dumper_213 = new("./depth213.csv");
    cstatus_csv_dumper_213 = new("./chan_status213.csv");
    fifo_monitor_213 = new(fifo_csv_dumper_213,fifo_intf_213,cstatus_csv_dumper_213);
    fifo_csv_dumper_214 = new("./depth214.csv");
    cstatus_csv_dumper_214 = new("./chan_status214.csv");
    fifo_monitor_214 = new(fifo_csv_dumper_214,fifo_intf_214,cstatus_csv_dumper_214);
    fifo_csv_dumper_215 = new("./depth215.csv");
    cstatus_csv_dumper_215 = new("./chan_status215.csv");
    fifo_monitor_215 = new(fifo_csv_dumper_215,fifo_intf_215,cstatus_csv_dumper_215);
    fifo_csv_dumper_216 = new("./depth216.csv");
    cstatus_csv_dumper_216 = new("./chan_status216.csv");
    fifo_monitor_216 = new(fifo_csv_dumper_216,fifo_intf_216,cstatus_csv_dumper_216);
    fifo_csv_dumper_217 = new("./depth217.csv");
    cstatus_csv_dumper_217 = new("./chan_status217.csv");
    fifo_monitor_217 = new(fifo_csv_dumper_217,fifo_intf_217,cstatus_csv_dumper_217);
    fifo_csv_dumper_218 = new("./depth218.csv");
    cstatus_csv_dumper_218 = new("./chan_status218.csv");
    fifo_monitor_218 = new(fifo_csv_dumper_218,fifo_intf_218,cstatus_csv_dumper_218);
    fifo_csv_dumper_219 = new("./depth219.csv");
    cstatus_csv_dumper_219 = new("./chan_status219.csv");
    fifo_monitor_219 = new(fifo_csv_dumper_219,fifo_intf_219,cstatus_csv_dumper_219);
    fifo_csv_dumper_220 = new("./depth220.csv");
    cstatus_csv_dumper_220 = new("./chan_status220.csv");
    fifo_monitor_220 = new(fifo_csv_dumper_220,fifo_intf_220,cstatus_csv_dumper_220);
    fifo_csv_dumper_221 = new("./depth221.csv");
    cstatus_csv_dumper_221 = new("./chan_status221.csv");
    fifo_monitor_221 = new(fifo_csv_dumper_221,fifo_intf_221,cstatus_csv_dumper_221);
    fifo_csv_dumper_222 = new("./depth222.csv");
    cstatus_csv_dumper_222 = new("./chan_status222.csv");
    fifo_monitor_222 = new(fifo_csv_dumper_222,fifo_intf_222,cstatus_csv_dumper_222);
    fifo_csv_dumper_223 = new("./depth223.csv");
    cstatus_csv_dumper_223 = new("./chan_status223.csv");
    fifo_monitor_223 = new(fifo_csv_dumper_223,fifo_intf_223,cstatus_csv_dumper_223);
    fifo_csv_dumper_224 = new("./depth224.csv");
    cstatus_csv_dumper_224 = new("./chan_status224.csv");
    fifo_monitor_224 = new(fifo_csv_dumper_224,fifo_intf_224,cstatus_csv_dumper_224);
    fifo_csv_dumper_225 = new("./depth225.csv");
    cstatus_csv_dumper_225 = new("./chan_status225.csv");
    fifo_monitor_225 = new(fifo_csv_dumper_225,fifo_intf_225,cstatus_csv_dumper_225);
    fifo_csv_dumper_226 = new("./depth226.csv");
    cstatus_csv_dumper_226 = new("./chan_status226.csv");
    fifo_monitor_226 = new(fifo_csv_dumper_226,fifo_intf_226,cstatus_csv_dumper_226);
    fifo_csv_dumper_227 = new("./depth227.csv");
    cstatus_csv_dumper_227 = new("./chan_status227.csv");
    fifo_monitor_227 = new(fifo_csv_dumper_227,fifo_intf_227,cstatus_csv_dumper_227);
    fifo_csv_dumper_228 = new("./depth228.csv");
    cstatus_csv_dumper_228 = new("./chan_status228.csv");
    fifo_monitor_228 = new(fifo_csv_dumper_228,fifo_intf_228,cstatus_csv_dumper_228);
    fifo_csv_dumper_229 = new("./depth229.csv");
    cstatus_csv_dumper_229 = new("./chan_status229.csv");
    fifo_monitor_229 = new(fifo_csv_dumper_229,fifo_intf_229,cstatus_csv_dumper_229);
    fifo_csv_dumper_230 = new("./depth230.csv");
    cstatus_csv_dumper_230 = new("./chan_status230.csv");
    fifo_monitor_230 = new(fifo_csv_dumper_230,fifo_intf_230,cstatus_csv_dumper_230);
    fifo_csv_dumper_231 = new("./depth231.csv");
    cstatus_csv_dumper_231 = new("./chan_status231.csv");
    fifo_monitor_231 = new(fifo_csv_dumper_231,fifo_intf_231,cstatus_csv_dumper_231);
    fifo_csv_dumper_232 = new("./depth232.csv");
    cstatus_csv_dumper_232 = new("./chan_status232.csv");
    fifo_monitor_232 = new(fifo_csv_dumper_232,fifo_intf_232,cstatus_csv_dumper_232);
    fifo_csv_dumper_233 = new("./depth233.csv");
    cstatus_csv_dumper_233 = new("./chan_status233.csv");
    fifo_monitor_233 = new(fifo_csv_dumper_233,fifo_intf_233,cstatus_csv_dumper_233);
    fifo_csv_dumper_234 = new("./depth234.csv");
    cstatus_csv_dumper_234 = new("./chan_status234.csv");
    fifo_monitor_234 = new(fifo_csv_dumper_234,fifo_intf_234,cstatus_csv_dumper_234);
    fifo_csv_dumper_235 = new("./depth235.csv");
    cstatus_csv_dumper_235 = new("./chan_status235.csv");
    fifo_monitor_235 = new(fifo_csv_dumper_235,fifo_intf_235,cstatus_csv_dumper_235);
    fifo_csv_dumper_236 = new("./depth236.csv");
    cstatus_csv_dumper_236 = new("./chan_status236.csv");
    fifo_monitor_236 = new(fifo_csv_dumper_236,fifo_intf_236,cstatus_csv_dumper_236);
    fifo_csv_dumper_237 = new("./depth237.csv");
    cstatus_csv_dumper_237 = new("./chan_status237.csv");
    fifo_monitor_237 = new(fifo_csv_dumper_237,fifo_intf_237,cstatus_csv_dumper_237);
    fifo_csv_dumper_238 = new("./depth238.csv");
    cstatus_csv_dumper_238 = new("./chan_status238.csv");
    fifo_monitor_238 = new(fifo_csv_dumper_238,fifo_intf_238,cstatus_csv_dumper_238);
    fifo_csv_dumper_239 = new("./depth239.csv");
    cstatus_csv_dumper_239 = new("./chan_status239.csv");
    fifo_monitor_239 = new(fifo_csv_dumper_239,fifo_intf_239,cstatus_csv_dumper_239);
    fifo_csv_dumper_240 = new("./depth240.csv");
    cstatus_csv_dumper_240 = new("./chan_status240.csv");
    fifo_monitor_240 = new(fifo_csv_dumper_240,fifo_intf_240,cstatus_csv_dumper_240);
    fifo_csv_dumper_241 = new("./depth241.csv");
    cstatus_csv_dumper_241 = new("./chan_status241.csv");
    fifo_monitor_241 = new(fifo_csv_dumper_241,fifo_intf_241,cstatus_csv_dumper_241);
    fifo_csv_dumper_242 = new("./depth242.csv");
    cstatus_csv_dumper_242 = new("./chan_status242.csv");
    fifo_monitor_242 = new(fifo_csv_dumper_242,fifo_intf_242,cstatus_csv_dumper_242);
    fifo_csv_dumper_243 = new("./depth243.csv");
    cstatus_csv_dumper_243 = new("./chan_status243.csv");
    fifo_monitor_243 = new(fifo_csv_dumper_243,fifo_intf_243,cstatus_csv_dumper_243);
    fifo_csv_dumper_244 = new("./depth244.csv");
    cstatus_csv_dumper_244 = new("./chan_status244.csv");
    fifo_monitor_244 = new(fifo_csv_dumper_244,fifo_intf_244,cstatus_csv_dumper_244);
    fifo_csv_dumper_245 = new("./depth245.csv");
    cstatus_csv_dumper_245 = new("./chan_status245.csv");
    fifo_monitor_245 = new(fifo_csv_dumper_245,fifo_intf_245,cstatus_csv_dumper_245);
    fifo_csv_dumper_246 = new("./depth246.csv");
    cstatus_csv_dumper_246 = new("./chan_status246.csv");
    fifo_monitor_246 = new(fifo_csv_dumper_246,fifo_intf_246,cstatus_csv_dumper_246);
    fifo_csv_dumper_247 = new("./depth247.csv");
    cstatus_csv_dumper_247 = new("./chan_status247.csv");
    fifo_monitor_247 = new(fifo_csv_dumper_247,fifo_intf_247,cstatus_csv_dumper_247);
    fifo_csv_dumper_248 = new("./depth248.csv");
    cstatus_csv_dumper_248 = new("./chan_status248.csv");
    fifo_monitor_248 = new(fifo_csv_dumper_248,fifo_intf_248,cstatus_csv_dumper_248);
    fifo_csv_dumper_249 = new("./depth249.csv");
    cstatus_csv_dumper_249 = new("./chan_status249.csv");
    fifo_monitor_249 = new(fifo_csv_dumper_249,fifo_intf_249,cstatus_csv_dumper_249);
    fifo_csv_dumper_250 = new("./depth250.csv");
    cstatus_csv_dumper_250 = new("./chan_status250.csv");
    fifo_monitor_250 = new(fifo_csv_dumper_250,fifo_intf_250,cstatus_csv_dumper_250);
    fifo_csv_dumper_251 = new("./depth251.csv");
    cstatus_csv_dumper_251 = new("./chan_status251.csv");
    fifo_monitor_251 = new(fifo_csv_dumper_251,fifo_intf_251,cstatus_csv_dumper_251);
    fifo_csv_dumper_252 = new("./depth252.csv");
    cstatus_csv_dumper_252 = new("./chan_status252.csv");
    fifo_monitor_252 = new(fifo_csv_dumper_252,fifo_intf_252,cstatus_csv_dumper_252);
    fifo_csv_dumper_253 = new("./depth253.csv");
    cstatus_csv_dumper_253 = new("./chan_status253.csv");
    fifo_monitor_253 = new(fifo_csv_dumper_253,fifo_intf_253,cstatus_csv_dumper_253);
    fifo_csv_dumper_254 = new("./depth254.csv");
    cstatus_csv_dumper_254 = new("./chan_status254.csv");
    fifo_monitor_254 = new(fifo_csv_dumper_254,fifo_intf_254,cstatus_csv_dumper_254);
    fifo_csv_dumper_255 = new("./depth255.csv");
    cstatus_csv_dumper_255 = new("./chan_status255.csv");
    fifo_monitor_255 = new(fifo_csv_dumper_255,fifo_intf_255,cstatus_csv_dumper_255);
    fifo_csv_dumper_256 = new("./depth256.csv");
    cstatus_csv_dumper_256 = new("./chan_status256.csv");
    fifo_monitor_256 = new(fifo_csv_dumper_256,fifo_intf_256,cstatus_csv_dumper_256);
    fifo_csv_dumper_257 = new("./depth257.csv");
    cstatus_csv_dumper_257 = new("./chan_status257.csv");
    fifo_monitor_257 = new(fifo_csv_dumper_257,fifo_intf_257,cstatus_csv_dumper_257);
    fifo_csv_dumper_258 = new("./depth258.csv");
    cstatus_csv_dumper_258 = new("./chan_status258.csv");
    fifo_monitor_258 = new(fifo_csv_dumper_258,fifo_intf_258,cstatus_csv_dumper_258);
    fifo_csv_dumper_259 = new("./depth259.csv");
    cstatus_csv_dumper_259 = new("./chan_status259.csv");
    fifo_monitor_259 = new(fifo_csv_dumper_259,fifo_intf_259,cstatus_csv_dumper_259);
    fifo_csv_dumper_260 = new("./depth260.csv");
    cstatus_csv_dumper_260 = new("./chan_status260.csv");
    fifo_monitor_260 = new(fifo_csv_dumper_260,fifo_intf_260,cstatus_csv_dumper_260);
    fifo_csv_dumper_261 = new("./depth261.csv");
    cstatus_csv_dumper_261 = new("./chan_status261.csv");
    fifo_monitor_261 = new(fifo_csv_dumper_261,fifo_intf_261,cstatus_csv_dumper_261);
    fifo_csv_dumper_262 = new("./depth262.csv");
    cstatus_csv_dumper_262 = new("./chan_status262.csv");
    fifo_monitor_262 = new(fifo_csv_dumper_262,fifo_intf_262,cstatus_csv_dumper_262);
    fifo_csv_dumper_263 = new("./depth263.csv");
    cstatus_csv_dumper_263 = new("./chan_status263.csv");
    fifo_monitor_263 = new(fifo_csv_dumper_263,fifo_intf_263,cstatus_csv_dumper_263);
    fifo_csv_dumper_264 = new("./depth264.csv");
    cstatus_csv_dumper_264 = new("./chan_status264.csv");
    fifo_monitor_264 = new(fifo_csv_dumper_264,fifo_intf_264,cstatus_csv_dumper_264);
    fifo_csv_dumper_265 = new("./depth265.csv");
    cstatus_csv_dumper_265 = new("./chan_status265.csv");
    fifo_monitor_265 = new(fifo_csv_dumper_265,fifo_intf_265,cstatus_csv_dumper_265);
    fifo_csv_dumper_266 = new("./depth266.csv");
    cstatus_csv_dumper_266 = new("./chan_status266.csv");
    fifo_monitor_266 = new(fifo_csv_dumper_266,fifo_intf_266,cstatus_csv_dumper_266);
    fifo_csv_dumper_267 = new("./depth267.csv");
    cstatus_csv_dumper_267 = new("./chan_status267.csv");
    fifo_monitor_267 = new(fifo_csv_dumper_267,fifo_intf_267,cstatus_csv_dumper_267);
    fifo_csv_dumper_268 = new("./depth268.csv");
    cstatus_csv_dumper_268 = new("./chan_status268.csv");
    fifo_monitor_268 = new(fifo_csv_dumper_268,fifo_intf_268,cstatus_csv_dumper_268);
    fifo_csv_dumper_269 = new("./depth269.csv");
    cstatus_csv_dumper_269 = new("./chan_status269.csv");
    fifo_monitor_269 = new(fifo_csv_dumper_269,fifo_intf_269,cstatus_csv_dumper_269);
    fifo_csv_dumper_270 = new("./depth270.csv");
    cstatus_csv_dumper_270 = new("./chan_status270.csv");
    fifo_monitor_270 = new(fifo_csv_dumper_270,fifo_intf_270,cstatus_csv_dumper_270);
    fifo_csv_dumper_271 = new("./depth271.csv");
    cstatus_csv_dumper_271 = new("./chan_status271.csv");
    fifo_monitor_271 = new(fifo_csv_dumper_271,fifo_intf_271,cstatus_csv_dumper_271);
    fifo_csv_dumper_272 = new("./depth272.csv");
    cstatus_csv_dumper_272 = new("./chan_status272.csv");
    fifo_monitor_272 = new(fifo_csv_dumper_272,fifo_intf_272,cstatus_csv_dumper_272);
    fifo_csv_dumper_273 = new("./depth273.csv");
    cstatus_csv_dumper_273 = new("./chan_status273.csv");
    fifo_monitor_273 = new(fifo_csv_dumper_273,fifo_intf_273,cstatus_csv_dumper_273);
    fifo_csv_dumper_274 = new("./depth274.csv");
    cstatus_csv_dumper_274 = new("./chan_status274.csv");
    fifo_monitor_274 = new(fifo_csv_dumper_274,fifo_intf_274,cstatus_csv_dumper_274);
    fifo_csv_dumper_275 = new("./depth275.csv");
    cstatus_csv_dumper_275 = new("./chan_status275.csv");
    fifo_monitor_275 = new(fifo_csv_dumper_275,fifo_intf_275,cstatus_csv_dumper_275);
    fifo_csv_dumper_276 = new("./depth276.csv");
    cstatus_csv_dumper_276 = new("./chan_status276.csv");
    fifo_monitor_276 = new(fifo_csv_dumper_276,fifo_intf_276,cstatus_csv_dumper_276);
    fifo_csv_dumper_277 = new("./depth277.csv");
    cstatus_csv_dumper_277 = new("./chan_status277.csv");
    fifo_monitor_277 = new(fifo_csv_dumper_277,fifo_intf_277,cstatus_csv_dumper_277);
    fifo_csv_dumper_278 = new("./depth278.csv");
    cstatus_csv_dumper_278 = new("./chan_status278.csv");
    fifo_monitor_278 = new(fifo_csv_dumper_278,fifo_intf_278,cstatus_csv_dumper_278);
    fifo_csv_dumper_279 = new("./depth279.csv");
    cstatus_csv_dumper_279 = new("./chan_status279.csv");
    fifo_monitor_279 = new(fifo_csv_dumper_279,fifo_intf_279,cstatus_csv_dumper_279);
    fifo_csv_dumper_280 = new("./depth280.csv");
    cstatus_csv_dumper_280 = new("./chan_status280.csv");
    fifo_monitor_280 = new(fifo_csv_dumper_280,fifo_intf_280,cstatus_csv_dumper_280);
    fifo_csv_dumper_281 = new("./depth281.csv");
    cstatus_csv_dumper_281 = new("./chan_status281.csv");
    fifo_monitor_281 = new(fifo_csv_dumper_281,fifo_intf_281,cstatus_csv_dumper_281);
    fifo_csv_dumper_282 = new("./depth282.csv");
    cstatus_csv_dumper_282 = new("./chan_status282.csv");
    fifo_monitor_282 = new(fifo_csv_dumper_282,fifo_intf_282,cstatus_csv_dumper_282);
    fifo_csv_dumper_283 = new("./depth283.csv");
    cstatus_csv_dumper_283 = new("./chan_status283.csv");
    fifo_monitor_283 = new(fifo_csv_dumper_283,fifo_intf_283,cstatus_csv_dumper_283);
    fifo_csv_dumper_284 = new("./depth284.csv");
    cstatus_csv_dumper_284 = new("./chan_status284.csv");
    fifo_monitor_284 = new(fifo_csv_dumper_284,fifo_intf_284,cstatus_csv_dumper_284);
    fifo_csv_dumper_285 = new("./depth285.csv");
    cstatus_csv_dumper_285 = new("./chan_status285.csv");
    fifo_monitor_285 = new(fifo_csv_dumper_285,fifo_intf_285,cstatus_csv_dumper_285);
    fifo_csv_dumper_286 = new("./depth286.csv");
    cstatus_csv_dumper_286 = new("./chan_status286.csv");
    fifo_monitor_286 = new(fifo_csv_dumper_286,fifo_intf_286,cstatus_csv_dumper_286);
    fifo_csv_dumper_287 = new("./depth287.csv");
    cstatus_csv_dumper_287 = new("./chan_status287.csv");
    fifo_monitor_287 = new(fifo_csv_dumper_287,fifo_intf_287,cstatus_csv_dumper_287);
    fifo_csv_dumper_288 = new("./depth288.csv");
    cstatus_csv_dumper_288 = new("./chan_status288.csv");
    fifo_monitor_288 = new(fifo_csv_dumper_288,fifo_intf_288,cstatus_csv_dumper_288);
    fifo_csv_dumper_289 = new("./depth289.csv");
    cstatus_csv_dumper_289 = new("./chan_status289.csv");
    fifo_monitor_289 = new(fifo_csv_dumper_289,fifo_intf_289,cstatus_csv_dumper_289);
    fifo_csv_dumper_290 = new("./depth290.csv");
    cstatus_csv_dumper_290 = new("./chan_status290.csv");
    fifo_monitor_290 = new(fifo_csv_dumper_290,fifo_intf_290,cstatus_csv_dumper_290);
    fifo_csv_dumper_291 = new("./depth291.csv");
    cstatus_csv_dumper_291 = new("./chan_status291.csv");
    fifo_monitor_291 = new(fifo_csv_dumper_291,fifo_intf_291,cstatus_csv_dumper_291);
    fifo_csv_dumper_292 = new("./depth292.csv");
    cstatus_csv_dumper_292 = new("./chan_status292.csv");
    fifo_monitor_292 = new(fifo_csv_dumper_292,fifo_intf_292,cstatus_csv_dumper_292);
    fifo_csv_dumper_293 = new("./depth293.csv");
    cstatus_csv_dumper_293 = new("./chan_status293.csv");
    fifo_monitor_293 = new(fifo_csv_dumper_293,fifo_intf_293,cstatus_csv_dumper_293);
    fifo_csv_dumper_294 = new("./depth294.csv");
    cstatus_csv_dumper_294 = new("./chan_status294.csv");
    fifo_monitor_294 = new(fifo_csv_dumper_294,fifo_intf_294,cstatus_csv_dumper_294);
    fifo_csv_dumper_295 = new("./depth295.csv");
    cstatus_csv_dumper_295 = new("./chan_status295.csv");
    fifo_monitor_295 = new(fifo_csv_dumper_295,fifo_intf_295,cstatus_csv_dumper_295);
    fifo_csv_dumper_296 = new("./depth296.csv");
    cstatus_csv_dumper_296 = new("./chan_status296.csv");
    fifo_monitor_296 = new(fifo_csv_dumper_296,fifo_intf_296,cstatus_csv_dumper_296);
    fifo_csv_dumper_297 = new("./depth297.csv");
    cstatus_csv_dumper_297 = new("./chan_status297.csv");
    fifo_monitor_297 = new(fifo_csv_dumper_297,fifo_intf_297,cstatus_csv_dumper_297);
    fifo_csv_dumper_298 = new("./depth298.csv");
    cstatus_csv_dumper_298 = new("./chan_status298.csv");
    fifo_monitor_298 = new(fifo_csv_dumper_298,fifo_intf_298,cstatus_csv_dumper_298);
    fifo_csv_dumper_299 = new("./depth299.csv");
    cstatus_csv_dumper_299 = new("./chan_status299.csv");
    fifo_monitor_299 = new(fifo_csv_dumper_299,fifo_intf_299,cstatus_csv_dumper_299);
    fifo_csv_dumper_300 = new("./depth300.csv");
    cstatus_csv_dumper_300 = new("./chan_status300.csv");
    fifo_monitor_300 = new(fifo_csv_dumper_300,fifo_intf_300,cstatus_csv_dumper_300);
    fifo_csv_dumper_301 = new("./depth301.csv");
    cstatus_csv_dumper_301 = new("./chan_status301.csv");
    fifo_monitor_301 = new(fifo_csv_dumper_301,fifo_intf_301,cstatus_csv_dumper_301);
    fifo_csv_dumper_302 = new("./depth302.csv");
    cstatus_csv_dumper_302 = new("./chan_status302.csv");
    fifo_monitor_302 = new(fifo_csv_dumper_302,fifo_intf_302,cstatus_csv_dumper_302);
    fifo_csv_dumper_303 = new("./depth303.csv");
    cstatus_csv_dumper_303 = new("./chan_status303.csv");
    fifo_monitor_303 = new(fifo_csv_dumper_303,fifo_intf_303,cstatus_csv_dumper_303);
    fifo_csv_dumper_304 = new("./depth304.csv");
    cstatus_csv_dumper_304 = new("./chan_status304.csv");
    fifo_monitor_304 = new(fifo_csv_dumper_304,fifo_intf_304,cstatus_csv_dumper_304);
    fifo_csv_dumper_305 = new("./depth305.csv");
    cstatus_csv_dumper_305 = new("./chan_status305.csv");
    fifo_monitor_305 = new(fifo_csv_dumper_305,fifo_intf_305,cstatus_csv_dumper_305);
    fifo_csv_dumper_306 = new("./depth306.csv");
    cstatus_csv_dumper_306 = new("./chan_status306.csv");
    fifo_monitor_306 = new(fifo_csv_dumper_306,fifo_intf_306,cstatus_csv_dumper_306);
    fifo_csv_dumper_307 = new("./depth307.csv");
    cstatus_csv_dumper_307 = new("./chan_status307.csv");
    fifo_monitor_307 = new(fifo_csv_dumper_307,fifo_intf_307,cstatus_csv_dumper_307);
    fifo_csv_dumper_308 = new("./depth308.csv");
    cstatus_csv_dumper_308 = new("./chan_status308.csv");
    fifo_monitor_308 = new(fifo_csv_dumper_308,fifo_intf_308,cstatus_csv_dumper_308);
    fifo_csv_dumper_309 = new("./depth309.csv");
    cstatus_csv_dumper_309 = new("./chan_status309.csv");
    fifo_monitor_309 = new(fifo_csv_dumper_309,fifo_intf_309,cstatus_csv_dumper_309);
    fifo_csv_dumper_310 = new("./depth310.csv");
    cstatus_csv_dumper_310 = new("./chan_status310.csv");
    fifo_monitor_310 = new(fifo_csv_dumper_310,fifo_intf_310,cstatus_csv_dumper_310);
    fifo_csv_dumper_311 = new("./depth311.csv");
    cstatus_csv_dumper_311 = new("./chan_status311.csv");
    fifo_monitor_311 = new(fifo_csv_dumper_311,fifo_intf_311,cstatus_csv_dumper_311);
    fifo_csv_dumper_312 = new("./depth312.csv");
    cstatus_csv_dumper_312 = new("./chan_status312.csv");
    fifo_monitor_312 = new(fifo_csv_dumper_312,fifo_intf_312,cstatus_csv_dumper_312);
    fifo_csv_dumper_313 = new("./depth313.csv");
    cstatus_csv_dumper_313 = new("./chan_status313.csv");
    fifo_monitor_313 = new(fifo_csv_dumper_313,fifo_intf_313,cstatus_csv_dumper_313);
    fifo_csv_dumper_314 = new("./depth314.csv");
    cstatus_csv_dumper_314 = new("./chan_status314.csv");
    fifo_monitor_314 = new(fifo_csv_dumper_314,fifo_intf_314,cstatus_csv_dumper_314);
    fifo_csv_dumper_315 = new("./depth315.csv");
    cstatus_csv_dumper_315 = new("./chan_status315.csv");
    fifo_monitor_315 = new(fifo_csv_dumper_315,fifo_intf_315,cstatus_csv_dumper_315);
    fifo_csv_dumper_316 = new("./depth316.csv");
    cstatus_csv_dumper_316 = new("./chan_status316.csv");
    fifo_monitor_316 = new(fifo_csv_dumper_316,fifo_intf_316,cstatus_csv_dumper_316);
    fifo_csv_dumper_317 = new("./depth317.csv");
    cstatus_csv_dumper_317 = new("./chan_status317.csv");
    fifo_monitor_317 = new(fifo_csv_dumper_317,fifo_intf_317,cstatus_csv_dumper_317);
    fifo_csv_dumper_318 = new("./depth318.csv");
    cstatus_csv_dumper_318 = new("./chan_status318.csv");
    fifo_monitor_318 = new(fifo_csv_dumper_318,fifo_intf_318,cstatus_csv_dumper_318);
    fifo_csv_dumper_319 = new("./depth319.csv");
    cstatus_csv_dumper_319 = new("./chan_status319.csv");
    fifo_monitor_319 = new(fifo_csv_dumper_319,fifo_intf_319,cstatus_csv_dumper_319);
    fifo_csv_dumper_320 = new("./depth320.csv");
    cstatus_csv_dumper_320 = new("./chan_status320.csv");
    fifo_monitor_320 = new(fifo_csv_dumper_320,fifo_intf_320,cstatus_csv_dumper_320);
    fifo_csv_dumper_321 = new("./depth321.csv");
    cstatus_csv_dumper_321 = new("./chan_status321.csv");
    fifo_monitor_321 = new(fifo_csv_dumper_321,fifo_intf_321,cstatus_csv_dumper_321);
    fifo_csv_dumper_322 = new("./depth322.csv");
    cstatus_csv_dumper_322 = new("./chan_status322.csv");
    fifo_monitor_322 = new(fifo_csv_dumper_322,fifo_intf_322,cstatus_csv_dumper_322);
    fifo_csv_dumper_323 = new("./depth323.csv");
    cstatus_csv_dumper_323 = new("./chan_status323.csv");
    fifo_monitor_323 = new(fifo_csv_dumper_323,fifo_intf_323,cstatus_csv_dumper_323);
    fifo_csv_dumper_324 = new("./depth324.csv");
    cstatus_csv_dumper_324 = new("./chan_status324.csv");
    fifo_monitor_324 = new(fifo_csv_dumper_324,fifo_intf_324,cstatus_csv_dumper_324);
    fifo_csv_dumper_325 = new("./depth325.csv");
    cstatus_csv_dumper_325 = new("./chan_status325.csv");
    fifo_monitor_325 = new(fifo_csv_dumper_325,fifo_intf_325,cstatus_csv_dumper_325);
    fifo_csv_dumper_326 = new("./depth326.csv");
    cstatus_csv_dumper_326 = new("./chan_status326.csv");
    fifo_monitor_326 = new(fifo_csv_dumper_326,fifo_intf_326,cstatus_csv_dumper_326);
    fifo_csv_dumper_327 = new("./depth327.csv");
    cstatus_csv_dumper_327 = new("./chan_status327.csv");
    fifo_monitor_327 = new(fifo_csv_dumper_327,fifo_intf_327,cstatus_csv_dumper_327);
    fifo_csv_dumper_328 = new("./depth328.csv");
    cstatus_csv_dumper_328 = new("./chan_status328.csv");
    fifo_monitor_328 = new(fifo_csv_dumper_328,fifo_intf_328,cstatus_csv_dumper_328);
    fifo_csv_dumper_329 = new("./depth329.csv");
    cstatus_csv_dumper_329 = new("./chan_status329.csv");
    fifo_monitor_329 = new(fifo_csv_dumper_329,fifo_intf_329,cstatus_csv_dumper_329);
    fifo_csv_dumper_330 = new("./depth330.csv");
    cstatus_csv_dumper_330 = new("./chan_status330.csv");
    fifo_monitor_330 = new(fifo_csv_dumper_330,fifo_intf_330,cstatus_csv_dumper_330);
    fifo_csv_dumper_331 = new("./depth331.csv");
    cstatus_csv_dumper_331 = new("./chan_status331.csv");
    fifo_monitor_331 = new(fifo_csv_dumper_331,fifo_intf_331,cstatus_csv_dumper_331);
    fifo_csv_dumper_332 = new("./depth332.csv");
    cstatus_csv_dumper_332 = new("./chan_status332.csv");
    fifo_monitor_332 = new(fifo_csv_dumper_332,fifo_intf_332,cstatus_csv_dumper_332);
    fifo_csv_dumper_333 = new("./depth333.csv");
    cstatus_csv_dumper_333 = new("./chan_status333.csv");
    fifo_monitor_333 = new(fifo_csv_dumper_333,fifo_intf_333,cstatus_csv_dumper_333);
    fifo_csv_dumper_334 = new("./depth334.csv");
    cstatus_csv_dumper_334 = new("./chan_status334.csv");
    fifo_monitor_334 = new(fifo_csv_dumper_334,fifo_intf_334,cstatus_csv_dumper_334);
    fifo_csv_dumper_335 = new("./depth335.csv");
    cstatus_csv_dumper_335 = new("./chan_status335.csv");
    fifo_monitor_335 = new(fifo_csv_dumper_335,fifo_intf_335,cstatus_csv_dumper_335);
    fifo_csv_dumper_336 = new("./depth336.csv");
    cstatus_csv_dumper_336 = new("./chan_status336.csv");
    fifo_monitor_336 = new(fifo_csv_dumper_336,fifo_intf_336,cstatus_csv_dumper_336);
    fifo_csv_dumper_337 = new("./depth337.csv");
    cstatus_csv_dumper_337 = new("./chan_status337.csv");
    fifo_monitor_337 = new(fifo_csv_dumper_337,fifo_intf_337,cstatus_csv_dumper_337);
    fifo_csv_dumper_338 = new("./depth338.csv");
    cstatus_csv_dumper_338 = new("./chan_status338.csv");
    fifo_monitor_338 = new(fifo_csv_dumper_338,fifo_intf_338,cstatus_csv_dumper_338);
    fifo_csv_dumper_339 = new("./depth339.csv");
    cstatus_csv_dumper_339 = new("./chan_status339.csv");
    fifo_monitor_339 = new(fifo_csv_dumper_339,fifo_intf_339,cstatus_csv_dumper_339);
    fifo_csv_dumper_340 = new("./depth340.csv");
    cstatus_csv_dumper_340 = new("./chan_status340.csv");
    fifo_monitor_340 = new(fifo_csv_dumper_340,fifo_intf_340,cstatus_csv_dumper_340);
    fifo_csv_dumper_341 = new("./depth341.csv");
    cstatus_csv_dumper_341 = new("./chan_status341.csv");
    fifo_monitor_341 = new(fifo_csv_dumper_341,fifo_intf_341,cstatus_csv_dumper_341);
    fifo_csv_dumper_342 = new("./depth342.csv");
    cstatus_csv_dumper_342 = new("./chan_status342.csv");
    fifo_monitor_342 = new(fifo_csv_dumper_342,fifo_intf_342,cstatus_csv_dumper_342);
    fifo_csv_dumper_343 = new("./depth343.csv");
    cstatus_csv_dumper_343 = new("./chan_status343.csv");
    fifo_monitor_343 = new(fifo_csv_dumper_343,fifo_intf_343,cstatus_csv_dumper_343);
    fifo_csv_dumper_344 = new("./depth344.csv");
    cstatus_csv_dumper_344 = new("./chan_status344.csv");
    fifo_monitor_344 = new(fifo_csv_dumper_344,fifo_intf_344,cstatus_csv_dumper_344);
    fifo_csv_dumper_345 = new("./depth345.csv");
    cstatus_csv_dumper_345 = new("./chan_status345.csv");
    fifo_monitor_345 = new(fifo_csv_dumper_345,fifo_intf_345,cstatus_csv_dumper_345);
    fifo_csv_dumper_346 = new("./depth346.csv");
    cstatus_csv_dumper_346 = new("./chan_status346.csv");
    fifo_monitor_346 = new(fifo_csv_dumper_346,fifo_intf_346,cstatus_csv_dumper_346);
    fifo_csv_dumper_347 = new("./depth347.csv");
    cstatus_csv_dumper_347 = new("./chan_status347.csv");
    fifo_monitor_347 = new(fifo_csv_dumper_347,fifo_intf_347,cstatus_csv_dumper_347);
    fifo_csv_dumper_348 = new("./depth348.csv");
    cstatus_csv_dumper_348 = new("./chan_status348.csv");
    fifo_monitor_348 = new(fifo_csv_dumper_348,fifo_intf_348,cstatus_csv_dumper_348);
    fifo_csv_dumper_349 = new("./depth349.csv");
    cstatus_csv_dumper_349 = new("./chan_status349.csv");
    fifo_monitor_349 = new(fifo_csv_dumper_349,fifo_intf_349,cstatus_csv_dumper_349);
    fifo_csv_dumper_350 = new("./depth350.csv");
    cstatus_csv_dumper_350 = new("./chan_status350.csv");
    fifo_monitor_350 = new(fifo_csv_dumper_350,fifo_intf_350,cstatus_csv_dumper_350);
    fifo_csv_dumper_351 = new("./depth351.csv");
    cstatus_csv_dumper_351 = new("./chan_status351.csv");
    fifo_monitor_351 = new(fifo_csv_dumper_351,fifo_intf_351,cstatus_csv_dumper_351);
    fifo_csv_dumper_352 = new("./depth352.csv");
    cstatus_csv_dumper_352 = new("./chan_status352.csv");
    fifo_monitor_352 = new(fifo_csv_dumper_352,fifo_intf_352,cstatus_csv_dumper_352);
    fifo_csv_dumper_353 = new("./depth353.csv");
    cstatus_csv_dumper_353 = new("./chan_status353.csv");
    fifo_monitor_353 = new(fifo_csv_dumper_353,fifo_intf_353,cstatus_csv_dumper_353);
    fifo_csv_dumper_354 = new("./depth354.csv");
    cstatus_csv_dumper_354 = new("./chan_status354.csv");
    fifo_monitor_354 = new(fifo_csv_dumper_354,fifo_intf_354,cstatus_csv_dumper_354);
    fifo_csv_dumper_355 = new("./depth355.csv");
    cstatus_csv_dumper_355 = new("./chan_status355.csv");
    fifo_monitor_355 = new(fifo_csv_dumper_355,fifo_intf_355,cstatus_csv_dumper_355);
    fifo_csv_dumper_356 = new("./depth356.csv");
    cstatus_csv_dumper_356 = new("./chan_status356.csv");
    fifo_monitor_356 = new(fifo_csv_dumper_356,fifo_intf_356,cstatus_csv_dumper_356);
    fifo_csv_dumper_357 = new("./depth357.csv");
    cstatus_csv_dumper_357 = new("./chan_status357.csv");
    fifo_monitor_357 = new(fifo_csv_dumper_357,fifo_intf_357,cstatus_csv_dumper_357);
    fifo_csv_dumper_358 = new("./depth358.csv");
    cstatus_csv_dumper_358 = new("./chan_status358.csv");
    fifo_monitor_358 = new(fifo_csv_dumper_358,fifo_intf_358,cstatus_csv_dumper_358);
    fifo_csv_dumper_359 = new("./depth359.csv");
    cstatus_csv_dumper_359 = new("./chan_status359.csv");
    fifo_monitor_359 = new(fifo_csv_dumper_359,fifo_intf_359,cstatus_csv_dumper_359);
    fifo_csv_dumper_360 = new("./depth360.csv");
    cstatus_csv_dumper_360 = new("./chan_status360.csv");
    fifo_monitor_360 = new(fifo_csv_dumper_360,fifo_intf_360,cstatus_csv_dumper_360);
    fifo_csv_dumper_361 = new("./depth361.csv");
    cstatus_csv_dumper_361 = new("./chan_status361.csv");
    fifo_monitor_361 = new(fifo_csv_dumper_361,fifo_intf_361,cstatus_csv_dumper_361);
    fifo_csv_dumper_362 = new("./depth362.csv");
    cstatus_csv_dumper_362 = new("./chan_status362.csv");
    fifo_monitor_362 = new(fifo_csv_dumper_362,fifo_intf_362,cstatus_csv_dumper_362);
    fifo_csv_dumper_363 = new("./depth363.csv");
    cstatus_csv_dumper_363 = new("./chan_status363.csv");
    fifo_monitor_363 = new(fifo_csv_dumper_363,fifo_intf_363,cstatus_csv_dumper_363);
    fifo_csv_dumper_364 = new("./depth364.csv");
    cstatus_csv_dumper_364 = new("./chan_status364.csv");
    fifo_monitor_364 = new(fifo_csv_dumper_364,fifo_intf_364,cstatus_csv_dumper_364);
    fifo_csv_dumper_365 = new("./depth365.csv");
    cstatus_csv_dumper_365 = new("./chan_status365.csv");
    fifo_monitor_365 = new(fifo_csv_dumper_365,fifo_intf_365,cstatus_csv_dumper_365);
    fifo_csv_dumper_366 = new("./depth366.csv");
    cstatus_csv_dumper_366 = new("./chan_status366.csv");
    fifo_monitor_366 = new(fifo_csv_dumper_366,fifo_intf_366,cstatus_csv_dumper_366);
    fifo_csv_dumper_367 = new("./depth367.csv");
    cstatus_csv_dumper_367 = new("./chan_status367.csv");
    fifo_monitor_367 = new(fifo_csv_dumper_367,fifo_intf_367,cstatus_csv_dumper_367);
    fifo_csv_dumper_368 = new("./depth368.csv");
    cstatus_csv_dumper_368 = new("./chan_status368.csv");
    fifo_monitor_368 = new(fifo_csv_dumper_368,fifo_intf_368,cstatus_csv_dumper_368);
    fifo_csv_dumper_369 = new("./depth369.csv");
    cstatus_csv_dumper_369 = new("./chan_status369.csv");
    fifo_monitor_369 = new(fifo_csv_dumper_369,fifo_intf_369,cstatus_csv_dumper_369);
    fifo_csv_dumper_370 = new("./depth370.csv");
    cstatus_csv_dumper_370 = new("./chan_status370.csv");
    fifo_monitor_370 = new(fifo_csv_dumper_370,fifo_intf_370,cstatus_csv_dumper_370);
    fifo_csv_dumper_371 = new("./depth371.csv");
    cstatus_csv_dumper_371 = new("./chan_status371.csv");
    fifo_monitor_371 = new(fifo_csv_dumper_371,fifo_intf_371,cstatus_csv_dumper_371);
    fifo_csv_dumper_372 = new("./depth372.csv");
    cstatus_csv_dumper_372 = new("./chan_status372.csv");
    fifo_monitor_372 = new(fifo_csv_dumper_372,fifo_intf_372,cstatus_csv_dumper_372);
    fifo_csv_dumper_373 = new("./depth373.csv");
    cstatus_csv_dumper_373 = new("./chan_status373.csv");
    fifo_monitor_373 = new(fifo_csv_dumper_373,fifo_intf_373,cstatus_csv_dumper_373);
    fifo_csv_dumper_374 = new("./depth374.csv");
    cstatus_csv_dumper_374 = new("./chan_status374.csv");
    fifo_monitor_374 = new(fifo_csv_dumper_374,fifo_intf_374,cstatus_csv_dumper_374);
    fifo_csv_dumper_375 = new("./depth375.csv");
    cstatus_csv_dumper_375 = new("./chan_status375.csv");
    fifo_monitor_375 = new(fifo_csv_dumper_375,fifo_intf_375,cstatus_csv_dumper_375);
    fifo_csv_dumper_376 = new("./depth376.csv");
    cstatus_csv_dumper_376 = new("./chan_status376.csv");
    fifo_monitor_376 = new(fifo_csv_dumper_376,fifo_intf_376,cstatus_csv_dumper_376);
    fifo_csv_dumper_377 = new("./depth377.csv");
    cstatus_csv_dumper_377 = new("./chan_status377.csv");
    fifo_monitor_377 = new(fifo_csv_dumper_377,fifo_intf_377,cstatus_csv_dumper_377);
    fifo_csv_dumper_378 = new("./depth378.csv");
    cstatus_csv_dumper_378 = new("./chan_status378.csv");
    fifo_monitor_378 = new(fifo_csv_dumper_378,fifo_intf_378,cstatus_csv_dumper_378);
    fifo_csv_dumper_379 = new("./depth379.csv");
    cstatus_csv_dumper_379 = new("./chan_status379.csv");
    fifo_monitor_379 = new(fifo_csv_dumper_379,fifo_intf_379,cstatus_csv_dumper_379);
    fifo_csv_dumper_380 = new("./depth380.csv");
    cstatus_csv_dumper_380 = new("./chan_status380.csv");
    fifo_monitor_380 = new(fifo_csv_dumper_380,fifo_intf_380,cstatus_csv_dumper_380);
    fifo_csv_dumper_381 = new("./depth381.csv");
    cstatus_csv_dumper_381 = new("./chan_status381.csv");
    fifo_monitor_381 = new(fifo_csv_dumper_381,fifo_intf_381,cstatus_csv_dumper_381);
    fifo_csv_dumper_382 = new("./depth382.csv");
    cstatus_csv_dumper_382 = new("./chan_status382.csv");
    fifo_monitor_382 = new(fifo_csv_dumper_382,fifo_intf_382,cstatus_csv_dumper_382);
    fifo_csv_dumper_383 = new("./depth383.csv");
    cstatus_csv_dumper_383 = new("./chan_status383.csv");
    fifo_monitor_383 = new(fifo_csv_dumper_383,fifo_intf_383,cstatus_csv_dumper_383);
    fifo_csv_dumper_384 = new("./depth384.csv");
    cstatus_csv_dumper_384 = new("./chan_status384.csv");
    fifo_monitor_384 = new(fifo_csv_dumper_384,fifo_intf_384,cstatus_csv_dumper_384);
    fifo_csv_dumper_385 = new("./depth385.csv");
    cstatus_csv_dumper_385 = new("./chan_status385.csv");
    fifo_monitor_385 = new(fifo_csv_dumper_385,fifo_intf_385,cstatus_csv_dumper_385);
    fifo_csv_dumper_386 = new("./depth386.csv");
    cstatus_csv_dumper_386 = new("./chan_status386.csv");
    fifo_monitor_386 = new(fifo_csv_dumper_386,fifo_intf_386,cstatus_csv_dumper_386);
    fifo_csv_dumper_387 = new("./depth387.csv");
    cstatus_csv_dumper_387 = new("./chan_status387.csv");
    fifo_monitor_387 = new(fifo_csv_dumper_387,fifo_intf_387,cstatus_csv_dumper_387);
    fifo_csv_dumper_388 = new("./depth388.csv");
    cstatus_csv_dumper_388 = new("./chan_status388.csv");
    fifo_monitor_388 = new(fifo_csv_dumper_388,fifo_intf_388,cstatus_csv_dumper_388);
    fifo_csv_dumper_389 = new("./depth389.csv");
    cstatus_csv_dumper_389 = new("./chan_status389.csv");
    fifo_monitor_389 = new(fifo_csv_dumper_389,fifo_intf_389,cstatus_csv_dumper_389);
    fifo_csv_dumper_390 = new("./depth390.csv");
    cstatus_csv_dumper_390 = new("./chan_status390.csv");
    fifo_monitor_390 = new(fifo_csv_dumper_390,fifo_intf_390,cstatus_csv_dumper_390);
    fifo_csv_dumper_391 = new("./depth391.csv");
    cstatus_csv_dumper_391 = new("./chan_status391.csv");
    fifo_monitor_391 = new(fifo_csv_dumper_391,fifo_intf_391,cstatus_csv_dumper_391);
    fifo_csv_dumper_392 = new("./depth392.csv");
    cstatus_csv_dumper_392 = new("./chan_status392.csv");
    fifo_monitor_392 = new(fifo_csv_dumper_392,fifo_intf_392,cstatus_csv_dumper_392);
    fifo_csv_dumper_393 = new("./depth393.csv");
    cstatus_csv_dumper_393 = new("./chan_status393.csv");
    fifo_monitor_393 = new(fifo_csv_dumper_393,fifo_intf_393,cstatus_csv_dumper_393);
    fifo_csv_dumper_394 = new("./depth394.csv");
    cstatus_csv_dumper_394 = new("./chan_status394.csv");
    fifo_monitor_394 = new(fifo_csv_dumper_394,fifo_intf_394,cstatus_csv_dumper_394);
    fifo_csv_dumper_395 = new("./depth395.csv");
    cstatus_csv_dumper_395 = new("./chan_status395.csv");
    fifo_monitor_395 = new(fifo_csv_dumper_395,fifo_intf_395,cstatus_csv_dumper_395);
    fifo_csv_dumper_396 = new("./depth396.csv");
    cstatus_csv_dumper_396 = new("./chan_status396.csv");
    fifo_monitor_396 = new(fifo_csv_dumper_396,fifo_intf_396,cstatus_csv_dumper_396);
    fifo_csv_dumper_397 = new("./depth397.csv");
    cstatus_csv_dumper_397 = new("./chan_status397.csv");
    fifo_monitor_397 = new(fifo_csv_dumper_397,fifo_intf_397,cstatus_csv_dumper_397);
    fifo_csv_dumper_398 = new("./depth398.csv");
    cstatus_csv_dumper_398 = new("./chan_status398.csv");
    fifo_monitor_398 = new(fifo_csv_dumper_398,fifo_intf_398,cstatus_csv_dumper_398);
    fifo_csv_dumper_399 = new("./depth399.csv");
    cstatus_csv_dumper_399 = new("./chan_status399.csv");
    fifo_monitor_399 = new(fifo_csv_dumper_399,fifo_intf_399,cstatus_csv_dumper_399);
    fifo_csv_dumper_400 = new("./depth400.csv");
    cstatus_csv_dumper_400 = new("./chan_status400.csv");
    fifo_monitor_400 = new(fifo_csv_dumper_400,fifo_intf_400,cstatus_csv_dumper_400);
    fifo_csv_dumper_401 = new("./depth401.csv");
    cstatus_csv_dumper_401 = new("./chan_status401.csv");
    fifo_monitor_401 = new(fifo_csv_dumper_401,fifo_intf_401,cstatus_csv_dumper_401);
    fifo_csv_dumper_402 = new("./depth402.csv");
    cstatus_csv_dumper_402 = new("./chan_status402.csv");
    fifo_monitor_402 = new(fifo_csv_dumper_402,fifo_intf_402,cstatus_csv_dumper_402);
    fifo_csv_dumper_403 = new("./depth403.csv");
    cstatus_csv_dumper_403 = new("./chan_status403.csv");
    fifo_monitor_403 = new(fifo_csv_dumper_403,fifo_intf_403,cstatus_csv_dumper_403);
    fifo_csv_dumper_404 = new("./depth404.csv");
    cstatus_csv_dumper_404 = new("./chan_status404.csv");
    fifo_monitor_404 = new(fifo_csv_dumper_404,fifo_intf_404,cstatus_csv_dumper_404);
    fifo_csv_dumper_405 = new("./depth405.csv");
    cstatus_csv_dumper_405 = new("./chan_status405.csv");
    fifo_monitor_405 = new(fifo_csv_dumper_405,fifo_intf_405,cstatus_csv_dumper_405);
    fifo_csv_dumper_406 = new("./depth406.csv");
    cstatus_csv_dumper_406 = new("./chan_status406.csv");
    fifo_monitor_406 = new(fifo_csv_dumper_406,fifo_intf_406,cstatus_csv_dumper_406);
    fifo_csv_dumper_407 = new("./depth407.csv");
    cstatus_csv_dumper_407 = new("./chan_status407.csv");
    fifo_monitor_407 = new(fifo_csv_dumper_407,fifo_intf_407,cstatus_csv_dumper_407);
    fifo_csv_dumper_408 = new("./depth408.csv");
    cstatus_csv_dumper_408 = new("./chan_status408.csv");
    fifo_monitor_408 = new(fifo_csv_dumper_408,fifo_intf_408,cstatus_csv_dumper_408);
    fifo_csv_dumper_409 = new("./depth409.csv");
    cstatus_csv_dumper_409 = new("./chan_status409.csv");
    fifo_monitor_409 = new(fifo_csv_dumper_409,fifo_intf_409,cstatus_csv_dumper_409);
    fifo_csv_dumper_410 = new("./depth410.csv");
    cstatus_csv_dumper_410 = new("./chan_status410.csv");
    fifo_monitor_410 = new(fifo_csv_dumper_410,fifo_intf_410,cstatus_csv_dumper_410);
    fifo_csv_dumper_411 = new("./depth411.csv");
    cstatus_csv_dumper_411 = new("./chan_status411.csv");
    fifo_monitor_411 = new(fifo_csv_dumper_411,fifo_intf_411,cstatus_csv_dumper_411);
    fifo_csv_dumper_412 = new("./depth412.csv");
    cstatus_csv_dumper_412 = new("./chan_status412.csv");
    fifo_monitor_412 = new(fifo_csv_dumper_412,fifo_intf_412,cstatus_csv_dumper_412);
    fifo_csv_dumper_413 = new("./depth413.csv");
    cstatus_csv_dumper_413 = new("./chan_status413.csv");
    fifo_monitor_413 = new(fifo_csv_dumper_413,fifo_intf_413,cstatus_csv_dumper_413);
    fifo_csv_dumper_414 = new("./depth414.csv");
    cstatus_csv_dumper_414 = new("./chan_status414.csv");
    fifo_monitor_414 = new(fifo_csv_dumper_414,fifo_intf_414,cstatus_csv_dumper_414);
    fifo_csv_dumper_415 = new("./depth415.csv");
    cstatus_csv_dumper_415 = new("./chan_status415.csv");
    fifo_monitor_415 = new(fifo_csv_dumper_415,fifo_intf_415,cstatus_csv_dumper_415);
    fifo_csv_dumper_416 = new("./depth416.csv");
    cstatus_csv_dumper_416 = new("./chan_status416.csv");
    fifo_monitor_416 = new(fifo_csv_dumper_416,fifo_intf_416,cstatus_csv_dumper_416);
    fifo_csv_dumper_417 = new("./depth417.csv");
    cstatus_csv_dumper_417 = new("./chan_status417.csv");
    fifo_monitor_417 = new(fifo_csv_dumper_417,fifo_intf_417,cstatus_csv_dumper_417);
    fifo_csv_dumper_418 = new("./depth418.csv");
    cstatus_csv_dumper_418 = new("./chan_status418.csv");
    fifo_monitor_418 = new(fifo_csv_dumper_418,fifo_intf_418,cstatus_csv_dumper_418);
    fifo_csv_dumper_419 = new("./depth419.csv");
    cstatus_csv_dumper_419 = new("./chan_status419.csv");
    fifo_monitor_419 = new(fifo_csv_dumper_419,fifo_intf_419,cstatus_csv_dumper_419);
    fifo_csv_dumper_420 = new("./depth420.csv");
    cstatus_csv_dumper_420 = new("./chan_status420.csv");
    fifo_monitor_420 = new(fifo_csv_dumper_420,fifo_intf_420,cstatus_csv_dumper_420);
    fifo_csv_dumper_421 = new("./depth421.csv");
    cstatus_csv_dumper_421 = new("./chan_status421.csv");
    fifo_monitor_421 = new(fifo_csv_dumper_421,fifo_intf_421,cstatus_csv_dumper_421);
    fifo_csv_dumper_422 = new("./depth422.csv");
    cstatus_csv_dumper_422 = new("./chan_status422.csv");
    fifo_monitor_422 = new(fifo_csv_dumper_422,fifo_intf_422,cstatus_csv_dumper_422);
    fifo_csv_dumper_423 = new("./depth423.csv");
    cstatus_csv_dumper_423 = new("./chan_status423.csv");
    fifo_monitor_423 = new(fifo_csv_dumper_423,fifo_intf_423,cstatus_csv_dumper_423);
    fifo_csv_dumper_424 = new("./depth424.csv");
    cstatus_csv_dumper_424 = new("./chan_status424.csv");
    fifo_monitor_424 = new(fifo_csv_dumper_424,fifo_intf_424,cstatus_csv_dumper_424);
    fifo_csv_dumper_425 = new("./depth425.csv");
    cstatus_csv_dumper_425 = new("./chan_status425.csv");
    fifo_monitor_425 = new(fifo_csv_dumper_425,fifo_intf_425,cstatus_csv_dumper_425);
    fifo_csv_dumper_426 = new("./depth426.csv");
    cstatus_csv_dumper_426 = new("./chan_status426.csv");
    fifo_monitor_426 = new(fifo_csv_dumper_426,fifo_intf_426,cstatus_csv_dumper_426);
    fifo_csv_dumper_427 = new("./depth427.csv");
    cstatus_csv_dumper_427 = new("./chan_status427.csv");
    fifo_monitor_427 = new(fifo_csv_dumper_427,fifo_intf_427,cstatus_csv_dumper_427);
    fifo_csv_dumper_428 = new("./depth428.csv");
    cstatus_csv_dumper_428 = new("./chan_status428.csv");
    fifo_monitor_428 = new(fifo_csv_dumper_428,fifo_intf_428,cstatus_csv_dumper_428);
    fifo_csv_dumper_429 = new("./depth429.csv");
    cstatus_csv_dumper_429 = new("./chan_status429.csv");
    fifo_monitor_429 = new(fifo_csv_dumper_429,fifo_intf_429,cstatus_csv_dumper_429);
    fifo_csv_dumper_430 = new("./depth430.csv");
    cstatus_csv_dumper_430 = new("./chan_status430.csv");
    fifo_monitor_430 = new(fifo_csv_dumper_430,fifo_intf_430,cstatus_csv_dumper_430);
    fifo_csv_dumper_431 = new("./depth431.csv");
    cstatus_csv_dumper_431 = new("./chan_status431.csv");
    fifo_monitor_431 = new(fifo_csv_dumper_431,fifo_intf_431,cstatus_csv_dumper_431);
    fifo_csv_dumper_432 = new("./depth432.csv");
    cstatus_csv_dumper_432 = new("./chan_status432.csv");
    fifo_monitor_432 = new(fifo_csv_dumper_432,fifo_intf_432,cstatus_csv_dumper_432);
    fifo_csv_dumper_433 = new("./depth433.csv");
    cstatus_csv_dumper_433 = new("./chan_status433.csv");
    fifo_monitor_433 = new(fifo_csv_dumper_433,fifo_intf_433,cstatus_csv_dumper_433);
    fifo_csv_dumper_434 = new("./depth434.csv");
    cstatus_csv_dumper_434 = new("./chan_status434.csv");
    fifo_monitor_434 = new(fifo_csv_dumper_434,fifo_intf_434,cstatus_csv_dumper_434);
    fifo_csv_dumper_435 = new("./depth435.csv");
    cstatus_csv_dumper_435 = new("./chan_status435.csv");
    fifo_monitor_435 = new(fifo_csv_dumper_435,fifo_intf_435,cstatus_csv_dumper_435);
    fifo_csv_dumper_436 = new("./depth436.csv");
    cstatus_csv_dumper_436 = new("./chan_status436.csv");
    fifo_monitor_436 = new(fifo_csv_dumper_436,fifo_intf_436,cstatus_csv_dumper_436);
    fifo_csv_dumper_437 = new("./depth437.csv");
    cstatus_csv_dumper_437 = new("./chan_status437.csv");
    fifo_monitor_437 = new(fifo_csv_dumper_437,fifo_intf_437,cstatus_csv_dumper_437);
    fifo_csv_dumper_438 = new("./depth438.csv");
    cstatus_csv_dumper_438 = new("./chan_status438.csv");
    fifo_monitor_438 = new(fifo_csv_dumper_438,fifo_intf_438,cstatus_csv_dumper_438);
    fifo_csv_dumper_439 = new("./depth439.csv");
    cstatus_csv_dumper_439 = new("./chan_status439.csv");
    fifo_monitor_439 = new(fifo_csv_dumper_439,fifo_intf_439,cstatus_csv_dumper_439);
    fifo_csv_dumper_440 = new("./depth440.csv");
    cstatus_csv_dumper_440 = new("./chan_status440.csv");
    fifo_monitor_440 = new(fifo_csv_dumper_440,fifo_intf_440,cstatus_csv_dumper_440);
    fifo_csv_dumper_441 = new("./depth441.csv");
    cstatus_csv_dumper_441 = new("./chan_status441.csv");
    fifo_monitor_441 = new(fifo_csv_dumper_441,fifo_intf_441,cstatus_csv_dumper_441);
    fifo_csv_dumper_442 = new("./depth442.csv");
    cstatus_csv_dumper_442 = new("./chan_status442.csv");
    fifo_monitor_442 = new(fifo_csv_dumper_442,fifo_intf_442,cstatus_csv_dumper_442);
    fifo_csv_dumper_443 = new("./depth443.csv");
    cstatus_csv_dumper_443 = new("./chan_status443.csv");
    fifo_monitor_443 = new(fifo_csv_dumper_443,fifo_intf_443,cstatus_csv_dumper_443);
    fifo_csv_dumper_444 = new("./depth444.csv");
    cstatus_csv_dumper_444 = new("./chan_status444.csv");
    fifo_monitor_444 = new(fifo_csv_dumper_444,fifo_intf_444,cstatus_csv_dumper_444);
    fifo_csv_dumper_445 = new("./depth445.csv");
    cstatus_csv_dumper_445 = new("./chan_status445.csv");
    fifo_monitor_445 = new(fifo_csv_dumper_445,fifo_intf_445,cstatus_csv_dumper_445);
    fifo_csv_dumper_446 = new("./depth446.csv");
    cstatus_csv_dumper_446 = new("./chan_status446.csv");
    fifo_monitor_446 = new(fifo_csv_dumper_446,fifo_intf_446,cstatus_csv_dumper_446);
    fifo_csv_dumper_447 = new("./depth447.csv");
    cstatus_csv_dumper_447 = new("./chan_status447.csv");
    fifo_monitor_447 = new(fifo_csv_dumper_447,fifo_intf_447,cstatus_csv_dumper_447);
    fifo_csv_dumper_448 = new("./depth448.csv");
    cstatus_csv_dumper_448 = new("./chan_status448.csv");
    fifo_monitor_448 = new(fifo_csv_dumper_448,fifo_intf_448,cstatus_csv_dumper_448);
    fifo_csv_dumper_449 = new("./depth449.csv");
    cstatus_csv_dumper_449 = new("./chan_status449.csv");
    fifo_monitor_449 = new(fifo_csv_dumper_449,fifo_intf_449,cstatus_csv_dumper_449);
    fifo_csv_dumper_450 = new("./depth450.csv");
    cstatus_csv_dumper_450 = new("./chan_status450.csv");
    fifo_monitor_450 = new(fifo_csv_dumper_450,fifo_intf_450,cstatus_csv_dumper_450);
    fifo_csv_dumper_451 = new("./depth451.csv");
    cstatus_csv_dumper_451 = new("./chan_status451.csv");
    fifo_monitor_451 = new(fifo_csv_dumper_451,fifo_intf_451,cstatus_csv_dumper_451);
    fifo_csv_dumper_452 = new("./depth452.csv");
    cstatus_csv_dumper_452 = new("./chan_status452.csv");
    fifo_monitor_452 = new(fifo_csv_dumper_452,fifo_intf_452,cstatus_csv_dumper_452);
    fifo_csv_dumper_453 = new("./depth453.csv");
    cstatus_csv_dumper_453 = new("./chan_status453.csv");
    fifo_monitor_453 = new(fifo_csv_dumper_453,fifo_intf_453,cstatus_csv_dumper_453);
    fifo_csv_dumper_454 = new("./depth454.csv");
    cstatus_csv_dumper_454 = new("./chan_status454.csv");
    fifo_monitor_454 = new(fifo_csv_dumper_454,fifo_intf_454,cstatus_csv_dumper_454);
    fifo_csv_dumper_455 = new("./depth455.csv");
    cstatus_csv_dumper_455 = new("./chan_status455.csv");
    fifo_monitor_455 = new(fifo_csv_dumper_455,fifo_intf_455,cstatus_csv_dumper_455);
    fifo_csv_dumper_456 = new("./depth456.csv");
    cstatus_csv_dumper_456 = new("./chan_status456.csv");
    fifo_monitor_456 = new(fifo_csv_dumper_456,fifo_intf_456,cstatus_csv_dumper_456);
    fifo_csv_dumper_457 = new("./depth457.csv");
    cstatus_csv_dumper_457 = new("./chan_status457.csv");
    fifo_monitor_457 = new(fifo_csv_dumper_457,fifo_intf_457,cstatus_csv_dumper_457);
    fifo_csv_dumper_458 = new("./depth458.csv");
    cstatus_csv_dumper_458 = new("./chan_status458.csv");
    fifo_monitor_458 = new(fifo_csv_dumper_458,fifo_intf_458,cstatus_csv_dumper_458);
    fifo_csv_dumper_459 = new("./depth459.csv");
    cstatus_csv_dumper_459 = new("./chan_status459.csv");
    fifo_monitor_459 = new(fifo_csv_dumper_459,fifo_intf_459,cstatus_csv_dumper_459);
    fifo_csv_dumper_460 = new("./depth460.csv");
    cstatus_csv_dumper_460 = new("./chan_status460.csv");
    fifo_monitor_460 = new(fifo_csv_dumper_460,fifo_intf_460,cstatus_csv_dumper_460);
    fifo_csv_dumper_461 = new("./depth461.csv");
    cstatus_csv_dumper_461 = new("./chan_status461.csv");
    fifo_monitor_461 = new(fifo_csv_dumper_461,fifo_intf_461,cstatus_csv_dumper_461);
    fifo_csv_dumper_462 = new("./depth462.csv");
    cstatus_csv_dumper_462 = new("./chan_status462.csv");
    fifo_monitor_462 = new(fifo_csv_dumper_462,fifo_intf_462,cstatus_csv_dumper_462);
    fifo_csv_dumper_463 = new("./depth463.csv");
    cstatus_csv_dumper_463 = new("./chan_status463.csv");
    fifo_monitor_463 = new(fifo_csv_dumper_463,fifo_intf_463,cstatus_csv_dumper_463);
    fifo_csv_dumper_464 = new("./depth464.csv");
    cstatus_csv_dumper_464 = new("./chan_status464.csv");
    fifo_monitor_464 = new(fifo_csv_dumper_464,fifo_intf_464,cstatus_csv_dumper_464);
    fifo_csv_dumper_465 = new("./depth465.csv");
    cstatus_csv_dumper_465 = new("./chan_status465.csv");
    fifo_monitor_465 = new(fifo_csv_dumper_465,fifo_intf_465,cstatus_csv_dumper_465);
    fifo_csv_dumper_466 = new("./depth466.csv");
    cstatus_csv_dumper_466 = new("./chan_status466.csv");
    fifo_monitor_466 = new(fifo_csv_dumper_466,fifo_intf_466,cstatus_csv_dumper_466);
    fifo_csv_dumper_467 = new("./depth467.csv");
    cstatus_csv_dumper_467 = new("./chan_status467.csv");
    fifo_monitor_467 = new(fifo_csv_dumper_467,fifo_intf_467,cstatus_csv_dumper_467);
    fifo_csv_dumper_468 = new("./depth468.csv");
    cstatus_csv_dumper_468 = new("./chan_status468.csv");
    fifo_monitor_468 = new(fifo_csv_dumper_468,fifo_intf_468,cstatus_csv_dumper_468);
    fifo_csv_dumper_469 = new("./depth469.csv");
    cstatus_csv_dumper_469 = new("./chan_status469.csv");
    fifo_monitor_469 = new(fifo_csv_dumper_469,fifo_intf_469,cstatus_csv_dumper_469);
    fifo_csv_dumper_470 = new("./depth470.csv");
    cstatus_csv_dumper_470 = new("./chan_status470.csv");
    fifo_monitor_470 = new(fifo_csv_dumper_470,fifo_intf_470,cstatus_csv_dumper_470);
    fifo_csv_dumper_471 = new("./depth471.csv");
    cstatus_csv_dumper_471 = new("./chan_status471.csv");
    fifo_monitor_471 = new(fifo_csv_dumper_471,fifo_intf_471,cstatus_csv_dumper_471);
    fifo_csv_dumper_472 = new("./depth472.csv");
    cstatus_csv_dumper_472 = new("./chan_status472.csv");
    fifo_monitor_472 = new(fifo_csv_dumper_472,fifo_intf_472,cstatus_csv_dumper_472);
    fifo_csv_dumper_473 = new("./depth473.csv");
    cstatus_csv_dumper_473 = new("./chan_status473.csv");
    fifo_monitor_473 = new(fifo_csv_dumper_473,fifo_intf_473,cstatus_csv_dumper_473);
    fifo_csv_dumper_474 = new("./depth474.csv");
    cstatus_csv_dumper_474 = new("./chan_status474.csv");
    fifo_monitor_474 = new(fifo_csv_dumper_474,fifo_intf_474,cstatus_csv_dumper_474);
    fifo_csv_dumper_475 = new("./depth475.csv");
    cstatus_csv_dumper_475 = new("./chan_status475.csv");
    fifo_monitor_475 = new(fifo_csv_dumper_475,fifo_intf_475,cstatus_csv_dumper_475);
    fifo_csv_dumper_476 = new("./depth476.csv");
    cstatus_csv_dumper_476 = new("./chan_status476.csv");
    fifo_monitor_476 = new(fifo_csv_dumper_476,fifo_intf_476,cstatus_csv_dumper_476);
    fifo_csv_dumper_477 = new("./depth477.csv");
    cstatus_csv_dumper_477 = new("./chan_status477.csv");
    fifo_monitor_477 = new(fifo_csv_dumper_477,fifo_intf_477,cstatus_csv_dumper_477);
    fifo_csv_dumper_478 = new("./depth478.csv");
    cstatus_csv_dumper_478 = new("./chan_status478.csv");
    fifo_monitor_478 = new(fifo_csv_dumper_478,fifo_intf_478,cstatus_csv_dumper_478);
    fifo_csv_dumper_479 = new("./depth479.csv");
    cstatus_csv_dumper_479 = new("./chan_status479.csv");
    fifo_monitor_479 = new(fifo_csv_dumper_479,fifo_intf_479,cstatus_csv_dumper_479);
    fifo_csv_dumper_480 = new("./depth480.csv");
    cstatus_csv_dumper_480 = new("./chan_status480.csv");
    fifo_monitor_480 = new(fifo_csv_dumper_480,fifo_intf_480,cstatus_csv_dumper_480);
    fifo_csv_dumper_481 = new("./depth481.csv");
    cstatus_csv_dumper_481 = new("./chan_status481.csv");
    fifo_monitor_481 = new(fifo_csv_dumper_481,fifo_intf_481,cstatus_csv_dumper_481);
    fifo_csv_dumper_482 = new("./depth482.csv");
    cstatus_csv_dumper_482 = new("./chan_status482.csv");
    fifo_monitor_482 = new(fifo_csv_dumper_482,fifo_intf_482,cstatus_csv_dumper_482);
    fifo_csv_dumper_483 = new("./depth483.csv");
    cstatus_csv_dumper_483 = new("./chan_status483.csv");
    fifo_monitor_483 = new(fifo_csv_dumper_483,fifo_intf_483,cstatus_csv_dumper_483);
    fifo_csv_dumper_484 = new("./depth484.csv");
    cstatus_csv_dumper_484 = new("./chan_status484.csv");
    fifo_monitor_484 = new(fifo_csv_dumper_484,fifo_intf_484,cstatus_csv_dumper_484);
    fifo_csv_dumper_485 = new("./depth485.csv");
    cstatus_csv_dumper_485 = new("./chan_status485.csv");
    fifo_monitor_485 = new(fifo_csv_dumper_485,fifo_intf_485,cstatus_csv_dumper_485);
    fifo_csv_dumper_486 = new("./depth486.csv");
    cstatus_csv_dumper_486 = new("./chan_status486.csv");
    fifo_monitor_486 = new(fifo_csv_dumper_486,fifo_intf_486,cstatus_csv_dumper_486);
    fifo_csv_dumper_487 = new("./depth487.csv");
    cstatus_csv_dumper_487 = new("./chan_status487.csv");
    fifo_monitor_487 = new(fifo_csv_dumper_487,fifo_intf_487,cstatus_csv_dumper_487);
    fifo_csv_dumper_488 = new("./depth488.csv");
    cstatus_csv_dumper_488 = new("./chan_status488.csv");
    fifo_monitor_488 = new(fifo_csv_dumper_488,fifo_intf_488,cstatus_csv_dumper_488);
    fifo_csv_dumper_489 = new("./depth489.csv");
    cstatus_csv_dumper_489 = new("./chan_status489.csv");
    fifo_monitor_489 = new(fifo_csv_dumper_489,fifo_intf_489,cstatus_csv_dumper_489);
    fifo_csv_dumper_490 = new("./depth490.csv");
    cstatus_csv_dumper_490 = new("./chan_status490.csv");
    fifo_monitor_490 = new(fifo_csv_dumper_490,fifo_intf_490,cstatus_csv_dumper_490);
    fifo_csv_dumper_491 = new("./depth491.csv");
    cstatus_csv_dumper_491 = new("./chan_status491.csv");
    fifo_monitor_491 = new(fifo_csv_dumper_491,fifo_intf_491,cstatus_csv_dumper_491);
    fifo_csv_dumper_492 = new("./depth492.csv");
    cstatus_csv_dumper_492 = new("./chan_status492.csv");
    fifo_monitor_492 = new(fifo_csv_dumper_492,fifo_intf_492,cstatus_csv_dumper_492);
    fifo_csv_dumper_493 = new("./depth493.csv");
    cstatus_csv_dumper_493 = new("./chan_status493.csv");
    fifo_monitor_493 = new(fifo_csv_dumper_493,fifo_intf_493,cstatus_csv_dumper_493);
    fifo_csv_dumper_494 = new("./depth494.csv");
    cstatus_csv_dumper_494 = new("./chan_status494.csv");
    fifo_monitor_494 = new(fifo_csv_dumper_494,fifo_intf_494,cstatus_csv_dumper_494);
    fifo_csv_dumper_495 = new("./depth495.csv");
    cstatus_csv_dumper_495 = new("./chan_status495.csv");
    fifo_monitor_495 = new(fifo_csv_dumper_495,fifo_intf_495,cstatus_csv_dumper_495);
    fifo_csv_dumper_496 = new("./depth496.csv");
    cstatus_csv_dumper_496 = new("./chan_status496.csv");
    fifo_monitor_496 = new(fifo_csv_dumper_496,fifo_intf_496,cstatus_csv_dumper_496);
    fifo_csv_dumper_497 = new("./depth497.csv");
    cstatus_csv_dumper_497 = new("./chan_status497.csv");
    fifo_monitor_497 = new(fifo_csv_dumper_497,fifo_intf_497,cstatus_csv_dumper_497);
    fifo_csv_dumper_498 = new("./depth498.csv");
    cstatus_csv_dumper_498 = new("./chan_status498.csv");
    fifo_monitor_498 = new(fifo_csv_dumper_498,fifo_intf_498,cstatus_csv_dumper_498);
    fifo_csv_dumper_499 = new("./depth499.csv");
    cstatus_csv_dumper_499 = new("./chan_status499.csv");
    fifo_monitor_499 = new(fifo_csv_dumper_499,fifo_intf_499,cstatus_csv_dumper_499);
    fifo_csv_dumper_500 = new("./depth500.csv");
    cstatus_csv_dumper_500 = new("./chan_status500.csv");
    fifo_monitor_500 = new(fifo_csv_dumper_500,fifo_intf_500,cstatus_csv_dumper_500);
    fifo_csv_dumper_501 = new("./depth501.csv");
    cstatus_csv_dumper_501 = new("./chan_status501.csv");
    fifo_monitor_501 = new(fifo_csv_dumper_501,fifo_intf_501,cstatus_csv_dumper_501);
    fifo_csv_dumper_502 = new("./depth502.csv");
    cstatus_csv_dumper_502 = new("./chan_status502.csv");
    fifo_monitor_502 = new(fifo_csv_dumper_502,fifo_intf_502,cstatus_csv_dumper_502);
    fifo_csv_dumper_503 = new("./depth503.csv");
    cstatus_csv_dumper_503 = new("./chan_status503.csv");
    fifo_monitor_503 = new(fifo_csv_dumper_503,fifo_intf_503,cstatus_csv_dumper_503);
    fifo_csv_dumper_504 = new("./depth504.csv");
    cstatus_csv_dumper_504 = new("./chan_status504.csv");
    fifo_monitor_504 = new(fifo_csv_dumper_504,fifo_intf_504,cstatus_csv_dumper_504);
    fifo_csv_dumper_505 = new("./depth505.csv");
    cstatus_csv_dumper_505 = new("./chan_status505.csv");
    fifo_monitor_505 = new(fifo_csv_dumper_505,fifo_intf_505,cstatus_csv_dumper_505);
    fifo_csv_dumper_506 = new("./depth506.csv");
    cstatus_csv_dumper_506 = new("./chan_status506.csv");
    fifo_monitor_506 = new(fifo_csv_dumper_506,fifo_intf_506,cstatus_csv_dumper_506);
    fifo_csv_dumper_507 = new("./depth507.csv");
    cstatus_csv_dumper_507 = new("./chan_status507.csv");
    fifo_monitor_507 = new(fifo_csv_dumper_507,fifo_intf_507,cstatus_csv_dumper_507);
    fifo_csv_dumper_508 = new("./depth508.csv");
    cstatus_csv_dumper_508 = new("./chan_status508.csv");
    fifo_monitor_508 = new(fifo_csv_dumper_508,fifo_intf_508,cstatus_csv_dumper_508);
    fifo_csv_dumper_509 = new("./depth509.csv");
    cstatus_csv_dumper_509 = new("./chan_status509.csv");
    fifo_monitor_509 = new(fifo_csv_dumper_509,fifo_intf_509,cstatus_csv_dumper_509);
    fifo_csv_dumper_510 = new("./depth510.csv");
    cstatus_csv_dumper_510 = new("./chan_status510.csv");
    fifo_monitor_510 = new(fifo_csv_dumper_510,fifo_intf_510,cstatus_csv_dumper_510);
    fifo_csv_dumper_511 = new("./depth511.csv");
    cstatus_csv_dumper_511 = new("./chan_status511.csv");
    fifo_monitor_511 = new(fifo_csv_dumper_511,fifo_intf_511,cstatus_csv_dumper_511);
    fifo_csv_dumper_512 = new("./depth512.csv");
    cstatus_csv_dumper_512 = new("./chan_status512.csv");
    fifo_monitor_512 = new(fifo_csv_dumper_512,fifo_intf_512,cstatus_csv_dumper_512);
    fifo_csv_dumper_513 = new("./depth513.csv");
    cstatus_csv_dumper_513 = new("./chan_status513.csv");
    fifo_monitor_513 = new(fifo_csv_dumper_513,fifo_intf_513,cstatus_csv_dumper_513);
    fifo_csv_dumper_514 = new("./depth514.csv");
    cstatus_csv_dumper_514 = new("./chan_status514.csv");
    fifo_monitor_514 = new(fifo_csv_dumper_514,fifo_intf_514,cstatus_csv_dumper_514);
    fifo_csv_dumper_515 = new("./depth515.csv");
    cstatus_csv_dumper_515 = new("./chan_status515.csv");
    fifo_monitor_515 = new(fifo_csv_dumper_515,fifo_intf_515,cstatus_csv_dumper_515);
    fifo_csv_dumper_516 = new("./depth516.csv");
    cstatus_csv_dumper_516 = new("./chan_status516.csv");
    fifo_monitor_516 = new(fifo_csv_dumper_516,fifo_intf_516,cstatus_csv_dumper_516);
    fifo_csv_dumper_517 = new("./depth517.csv");
    cstatus_csv_dumper_517 = new("./chan_status517.csv");
    fifo_monitor_517 = new(fifo_csv_dumper_517,fifo_intf_517,cstatus_csv_dumper_517);
    fifo_csv_dumper_518 = new("./depth518.csv");
    cstatus_csv_dumper_518 = new("./chan_status518.csv");
    fifo_monitor_518 = new(fifo_csv_dumper_518,fifo_intf_518,cstatus_csv_dumper_518);
    fifo_csv_dumper_519 = new("./depth519.csv");
    cstatus_csv_dumper_519 = new("./chan_status519.csv");
    fifo_monitor_519 = new(fifo_csv_dumper_519,fifo_intf_519,cstatus_csv_dumper_519);
    fifo_csv_dumper_520 = new("./depth520.csv");
    cstatus_csv_dumper_520 = new("./chan_status520.csv");
    fifo_monitor_520 = new(fifo_csv_dumper_520,fifo_intf_520,cstatus_csv_dumper_520);
    fifo_csv_dumper_521 = new("./depth521.csv");
    cstatus_csv_dumper_521 = new("./chan_status521.csv");
    fifo_monitor_521 = new(fifo_csv_dumper_521,fifo_intf_521,cstatus_csv_dumper_521);
    fifo_csv_dumper_522 = new("./depth522.csv");
    cstatus_csv_dumper_522 = new("./chan_status522.csv");
    fifo_monitor_522 = new(fifo_csv_dumper_522,fifo_intf_522,cstatus_csv_dumper_522);
    fifo_csv_dumper_523 = new("./depth523.csv");
    cstatus_csv_dumper_523 = new("./chan_status523.csv");
    fifo_monitor_523 = new(fifo_csv_dumper_523,fifo_intf_523,cstatus_csv_dumper_523);
    fifo_csv_dumper_524 = new("./depth524.csv");
    cstatus_csv_dumper_524 = new("./chan_status524.csv");
    fifo_monitor_524 = new(fifo_csv_dumper_524,fifo_intf_524,cstatus_csv_dumper_524);
    fifo_csv_dumper_525 = new("./depth525.csv");
    cstatus_csv_dumper_525 = new("./chan_status525.csv");
    fifo_monitor_525 = new(fifo_csv_dumper_525,fifo_intf_525,cstatus_csv_dumper_525);
    fifo_csv_dumper_526 = new("./depth526.csv");
    cstatus_csv_dumper_526 = new("./chan_status526.csv");
    fifo_monitor_526 = new(fifo_csv_dumper_526,fifo_intf_526,cstatus_csv_dumper_526);
    fifo_csv_dumper_527 = new("./depth527.csv");
    cstatus_csv_dumper_527 = new("./chan_status527.csv");
    fifo_monitor_527 = new(fifo_csv_dumper_527,fifo_intf_527,cstatus_csv_dumper_527);
    fifo_csv_dumper_528 = new("./depth528.csv");
    cstatus_csv_dumper_528 = new("./chan_status528.csv");
    fifo_monitor_528 = new(fifo_csv_dumper_528,fifo_intf_528,cstatus_csv_dumper_528);
    fifo_csv_dumper_529 = new("./depth529.csv");
    cstatus_csv_dumper_529 = new("./chan_status529.csv");
    fifo_monitor_529 = new(fifo_csv_dumper_529,fifo_intf_529,cstatus_csv_dumper_529);
    fifo_csv_dumper_530 = new("./depth530.csv");
    cstatus_csv_dumper_530 = new("./chan_status530.csv");
    fifo_monitor_530 = new(fifo_csv_dumper_530,fifo_intf_530,cstatus_csv_dumper_530);
    fifo_csv_dumper_531 = new("./depth531.csv");
    cstatus_csv_dumper_531 = new("./chan_status531.csv");
    fifo_monitor_531 = new(fifo_csv_dumper_531,fifo_intf_531,cstatus_csv_dumper_531);
    fifo_csv_dumper_532 = new("./depth532.csv");
    cstatus_csv_dumper_532 = new("./chan_status532.csv");
    fifo_monitor_532 = new(fifo_csv_dumper_532,fifo_intf_532,cstatus_csv_dumper_532);
    fifo_csv_dumper_533 = new("./depth533.csv");
    cstatus_csv_dumper_533 = new("./chan_status533.csv");
    fifo_monitor_533 = new(fifo_csv_dumper_533,fifo_intf_533,cstatus_csv_dumper_533);
    fifo_csv_dumper_534 = new("./depth534.csv");
    cstatus_csv_dumper_534 = new("./chan_status534.csv");
    fifo_monitor_534 = new(fifo_csv_dumper_534,fifo_intf_534,cstatus_csv_dumper_534);
    fifo_csv_dumper_535 = new("./depth535.csv");
    cstatus_csv_dumper_535 = new("./chan_status535.csv");
    fifo_monitor_535 = new(fifo_csv_dumper_535,fifo_intf_535,cstatus_csv_dumper_535);
    fifo_csv_dumper_536 = new("./depth536.csv");
    cstatus_csv_dumper_536 = new("./chan_status536.csv");
    fifo_monitor_536 = new(fifo_csv_dumper_536,fifo_intf_536,cstatus_csv_dumper_536);
    fifo_csv_dumper_537 = new("./depth537.csv");
    cstatus_csv_dumper_537 = new("./chan_status537.csv");
    fifo_monitor_537 = new(fifo_csv_dumper_537,fifo_intf_537,cstatus_csv_dumper_537);
    fifo_csv_dumper_538 = new("./depth538.csv");
    cstatus_csv_dumper_538 = new("./chan_status538.csv");
    fifo_monitor_538 = new(fifo_csv_dumper_538,fifo_intf_538,cstatus_csv_dumper_538);
    fifo_csv_dumper_539 = new("./depth539.csv");
    cstatus_csv_dumper_539 = new("./chan_status539.csv");
    fifo_monitor_539 = new(fifo_csv_dumper_539,fifo_intf_539,cstatus_csv_dumper_539);
    fifo_csv_dumper_540 = new("./depth540.csv");
    cstatus_csv_dumper_540 = new("./chan_status540.csv");
    fifo_monitor_540 = new(fifo_csv_dumper_540,fifo_intf_540,cstatus_csv_dumper_540);
    fifo_csv_dumper_541 = new("./depth541.csv");
    cstatus_csv_dumper_541 = new("./chan_status541.csv");
    fifo_monitor_541 = new(fifo_csv_dumper_541,fifo_intf_541,cstatus_csv_dumper_541);
    fifo_csv_dumper_542 = new("./depth542.csv");
    cstatus_csv_dumper_542 = new("./chan_status542.csv");
    fifo_monitor_542 = new(fifo_csv_dumper_542,fifo_intf_542,cstatus_csv_dumper_542);
    fifo_csv_dumper_543 = new("./depth543.csv");
    cstatus_csv_dumper_543 = new("./chan_status543.csv");
    fifo_monitor_543 = new(fifo_csv_dumper_543,fifo_intf_543,cstatus_csv_dumper_543);
    fifo_csv_dumper_544 = new("./depth544.csv");
    cstatus_csv_dumper_544 = new("./chan_status544.csv");
    fifo_monitor_544 = new(fifo_csv_dumper_544,fifo_intf_544,cstatus_csv_dumper_544);
    fifo_csv_dumper_545 = new("./depth545.csv");
    cstatus_csv_dumper_545 = new("./chan_status545.csv");
    fifo_monitor_545 = new(fifo_csv_dumper_545,fifo_intf_545,cstatus_csv_dumper_545);
    fifo_csv_dumper_546 = new("./depth546.csv");
    cstatus_csv_dumper_546 = new("./chan_status546.csv");
    fifo_monitor_546 = new(fifo_csv_dumper_546,fifo_intf_546,cstatus_csv_dumper_546);
    fifo_csv_dumper_547 = new("./depth547.csv");
    cstatus_csv_dumper_547 = new("./chan_status547.csv");
    fifo_monitor_547 = new(fifo_csv_dumper_547,fifo_intf_547,cstatus_csv_dumper_547);
    fifo_csv_dumper_548 = new("./depth548.csv");
    cstatus_csv_dumper_548 = new("./chan_status548.csv");
    fifo_monitor_548 = new(fifo_csv_dumper_548,fifo_intf_548,cstatus_csv_dumper_548);
    fifo_csv_dumper_549 = new("./depth549.csv");
    cstatus_csv_dumper_549 = new("./chan_status549.csv");
    fifo_monitor_549 = new(fifo_csv_dumper_549,fifo_intf_549,cstatus_csv_dumper_549);
    fifo_csv_dumper_550 = new("./depth550.csv");
    cstatus_csv_dumper_550 = new("./chan_status550.csv");
    fifo_monitor_550 = new(fifo_csv_dumper_550,fifo_intf_550,cstatus_csv_dumper_550);
    fifo_csv_dumper_551 = new("./depth551.csv");
    cstatus_csv_dumper_551 = new("./chan_status551.csv");
    fifo_monitor_551 = new(fifo_csv_dumper_551,fifo_intf_551,cstatus_csv_dumper_551);
    fifo_csv_dumper_552 = new("./depth552.csv");
    cstatus_csv_dumper_552 = new("./chan_status552.csv");
    fifo_monitor_552 = new(fifo_csv_dumper_552,fifo_intf_552,cstatus_csv_dumper_552);
    fifo_csv_dumper_553 = new("./depth553.csv");
    cstatus_csv_dumper_553 = new("./chan_status553.csv");
    fifo_monitor_553 = new(fifo_csv_dumper_553,fifo_intf_553,cstatus_csv_dumper_553);
    fifo_csv_dumper_554 = new("./depth554.csv");
    cstatus_csv_dumper_554 = new("./chan_status554.csv");
    fifo_monitor_554 = new(fifo_csv_dumper_554,fifo_intf_554,cstatus_csv_dumper_554);
    fifo_csv_dumper_555 = new("./depth555.csv");
    cstatus_csv_dumper_555 = new("./chan_status555.csv");
    fifo_monitor_555 = new(fifo_csv_dumper_555,fifo_intf_555,cstatus_csv_dumper_555);
    fifo_csv_dumper_556 = new("./depth556.csv");
    cstatus_csv_dumper_556 = new("./chan_status556.csv");
    fifo_monitor_556 = new(fifo_csv_dumper_556,fifo_intf_556,cstatus_csv_dumper_556);
    fifo_csv_dumper_557 = new("./depth557.csv");
    cstatus_csv_dumper_557 = new("./chan_status557.csv");
    fifo_monitor_557 = new(fifo_csv_dumper_557,fifo_intf_557,cstatus_csv_dumper_557);
    fifo_csv_dumper_558 = new("./depth558.csv");
    cstatus_csv_dumper_558 = new("./chan_status558.csv");
    fifo_monitor_558 = new(fifo_csv_dumper_558,fifo_intf_558,cstatus_csv_dumper_558);
    fifo_csv_dumper_559 = new("./depth559.csv");
    cstatus_csv_dumper_559 = new("./chan_status559.csv");
    fifo_monitor_559 = new(fifo_csv_dumper_559,fifo_intf_559,cstatus_csv_dumper_559);
    fifo_csv_dumper_560 = new("./depth560.csv");
    cstatus_csv_dumper_560 = new("./chan_status560.csv");
    fifo_monitor_560 = new(fifo_csv_dumper_560,fifo_intf_560,cstatus_csv_dumper_560);
    fifo_csv_dumper_561 = new("./depth561.csv");
    cstatus_csv_dumper_561 = new("./chan_status561.csv");
    fifo_monitor_561 = new(fifo_csv_dumper_561,fifo_intf_561,cstatus_csv_dumper_561);
    fifo_csv_dumper_562 = new("./depth562.csv");
    cstatus_csv_dumper_562 = new("./chan_status562.csv");
    fifo_monitor_562 = new(fifo_csv_dumper_562,fifo_intf_562,cstatus_csv_dumper_562);
    fifo_csv_dumper_563 = new("./depth563.csv");
    cstatus_csv_dumper_563 = new("./chan_status563.csv");
    fifo_monitor_563 = new(fifo_csv_dumper_563,fifo_intf_563,cstatus_csv_dumper_563);
    fifo_csv_dumper_564 = new("./depth564.csv");
    cstatus_csv_dumper_564 = new("./chan_status564.csv");
    fifo_monitor_564 = new(fifo_csv_dumper_564,fifo_intf_564,cstatus_csv_dumper_564);
    fifo_csv_dumper_565 = new("./depth565.csv");
    cstatus_csv_dumper_565 = new("./chan_status565.csv");
    fifo_monitor_565 = new(fifo_csv_dumper_565,fifo_intf_565,cstatus_csv_dumper_565);
    fifo_csv_dumper_566 = new("./depth566.csv");
    cstatus_csv_dumper_566 = new("./chan_status566.csv");
    fifo_monitor_566 = new(fifo_csv_dumper_566,fifo_intf_566,cstatus_csv_dumper_566);
    fifo_csv_dumper_567 = new("./depth567.csv");
    cstatus_csv_dumper_567 = new("./chan_status567.csv");
    fifo_monitor_567 = new(fifo_csv_dumper_567,fifo_intf_567,cstatus_csv_dumper_567);
    fifo_csv_dumper_568 = new("./depth568.csv");
    cstatus_csv_dumper_568 = new("./chan_status568.csv");
    fifo_monitor_568 = new(fifo_csv_dumper_568,fifo_intf_568,cstatus_csv_dumper_568);
    fifo_csv_dumper_569 = new("./depth569.csv");
    cstatus_csv_dumper_569 = new("./chan_status569.csv");
    fifo_monitor_569 = new(fifo_csv_dumper_569,fifo_intf_569,cstatus_csv_dumper_569);
    fifo_csv_dumper_570 = new("./depth570.csv");
    cstatus_csv_dumper_570 = new("./chan_status570.csv");
    fifo_monitor_570 = new(fifo_csv_dumper_570,fifo_intf_570,cstatus_csv_dumper_570);
    fifo_csv_dumper_571 = new("./depth571.csv");
    cstatus_csv_dumper_571 = new("./chan_status571.csv");
    fifo_monitor_571 = new(fifo_csv_dumper_571,fifo_intf_571,cstatus_csv_dumper_571);
    fifo_csv_dumper_572 = new("./depth572.csv");
    cstatus_csv_dumper_572 = new("./chan_status572.csv");
    fifo_monitor_572 = new(fifo_csv_dumper_572,fifo_intf_572,cstatus_csv_dumper_572);
    fifo_csv_dumper_573 = new("./depth573.csv");
    cstatus_csv_dumper_573 = new("./chan_status573.csv");
    fifo_monitor_573 = new(fifo_csv_dumper_573,fifo_intf_573,cstatus_csv_dumper_573);
    fifo_csv_dumper_574 = new("./depth574.csv");
    cstatus_csv_dumper_574 = new("./chan_status574.csv");
    fifo_monitor_574 = new(fifo_csv_dumper_574,fifo_intf_574,cstatus_csv_dumper_574);
    fifo_csv_dumper_575 = new("./depth575.csv");
    cstatus_csv_dumper_575 = new("./chan_status575.csv");
    fifo_monitor_575 = new(fifo_csv_dumper_575,fifo_intf_575,cstatus_csv_dumper_575);
    fifo_csv_dumper_576 = new("./depth576.csv");
    cstatus_csv_dumper_576 = new("./chan_status576.csv");
    fifo_monitor_576 = new(fifo_csv_dumper_576,fifo_intf_576,cstatus_csv_dumper_576);
    fifo_csv_dumper_577 = new("./depth577.csv");
    cstatus_csv_dumper_577 = new("./chan_status577.csv");
    fifo_monitor_577 = new(fifo_csv_dumper_577,fifo_intf_577,cstatus_csv_dumper_577);
    fifo_csv_dumper_578 = new("./depth578.csv");
    cstatus_csv_dumper_578 = new("./chan_status578.csv");
    fifo_monitor_578 = new(fifo_csv_dumper_578,fifo_intf_578,cstatus_csv_dumper_578);
    fifo_csv_dumper_579 = new("./depth579.csv");
    cstatus_csv_dumper_579 = new("./chan_status579.csv");
    fifo_monitor_579 = new(fifo_csv_dumper_579,fifo_intf_579,cstatus_csv_dumper_579);
    fifo_csv_dumper_580 = new("./depth580.csv");
    cstatus_csv_dumper_580 = new("./chan_status580.csv");
    fifo_monitor_580 = new(fifo_csv_dumper_580,fifo_intf_580,cstatus_csv_dumper_580);
    fifo_csv_dumper_581 = new("./depth581.csv");
    cstatus_csv_dumper_581 = new("./chan_status581.csv");
    fifo_monitor_581 = new(fifo_csv_dumper_581,fifo_intf_581,cstatus_csv_dumper_581);
    fifo_csv_dumper_582 = new("./depth582.csv");
    cstatus_csv_dumper_582 = new("./chan_status582.csv");
    fifo_monitor_582 = new(fifo_csv_dumper_582,fifo_intf_582,cstatus_csv_dumper_582);
    fifo_csv_dumper_583 = new("./depth583.csv");
    cstatus_csv_dumper_583 = new("./chan_status583.csv");
    fifo_monitor_583 = new(fifo_csv_dumper_583,fifo_intf_583,cstatus_csv_dumper_583);
    fifo_csv_dumper_584 = new("./depth584.csv");
    cstatus_csv_dumper_584 = new("./chan_status584.csv");
    fifo_monitor_584 = new(fifo_csv_dumper_584,fifo_intf_584,cstatus_csv_dumper_584);
    fifo_csv_dumper_585 = new("./depth585.csv");
    cstatus_csv_dumper_585 = new("./chan_status585.csv");
    fifo_monitor_585 = new(fifo_csv_dumper_585,fifo_intf_585,cstatus_csv_dumper_585);
    fifo_csv_dumper_586 = new("./depth586.csv");
    cstatus_csv_dumper_586 = new("./chan_status586.csv");
    fifo_monitor_586 = new(fifo_csv_dumper_586,fifo_intf_586,cstatus_csv_dumper_586);
    fifo_csv_dumper_587 = new("./depth587.csv");
    cstatus_csv_dumper_587 = new("./chan_status587.csv");
    fifo_monitor_587 = new(fifo_csv_dumper_587,fifo_intf_587,cstatus_csv_dumper_587);
    fifo_csv_dumper_588 = new("./depth588.csv");
    cstatus_csv_dumper_588 = new("./chan_status588.csv");
    fifo_monitor_588 = new(fifo_csv_dumper_588,fifo_intf_588,cstatus_csv_dumper_588);
    fifo_csv_dumper_589 = new("./depth589.csv");
    cstatus_csv_dumper_589 = new("./chan_status589.csv");
    fifo_monitor_589 = new(fifo_csv_dumper_589,fifo_intf_589,cstatus_csv_dumper_589);
    fifo_csv_dumper_590 = new("./depth590.csv");
    cstatus_csv_dumper_590 = new("./chan_status590.csv");
    fifo_monitor_590 = new(fifo_csv_dumper_590,fifo_intf_590,cstatus_csv_dumper_590);
    fifo_csv_dumper_591 = new("./depth591.csv");
    cstatus_csv_dumper_591 = new("./chan_status591.csv");
    fifo_monitor_591 = new(fifo_csv_dumper_591,fifo_intf_591,cstatus_csv_dumper_591);
    fifo_csv_dumper_592 = new("./depth592.csv");
    cstatus_csv_dumper_592 = new("./chan_status592.csv");
    fifo_monitor_592 = new(fifo_csv_dumper_592,fifo_intf_592,cstatus_csv_dumper_592);
    fifo_csv_dumper_593 = new("./depth593.csv");
    cstatus_csv_dumper_593 = new("./chan_status593.csv");
    fifo_monitor_593 = new(fifo_csv_dumper_593,fifo_intf_593,cstatus_csv_dumper_593);
    fifo_csv_dumper_594 = new("./depth594.csv");
    cstatus_csv_dumper_594 = new("./chan_status594.csv");
    fifo_monitor_594 = new(fifo_csv_dumper_594,fifo_intf_594,cstatus_csv_dumper_594);
    fifo_csv_dumper_595 = new("./depth595.csv");
    cstatus_csv_dumper_595 = new("./chan_status595.csv");
    fifo_monitor_595 = new(fifo_csv_dumper_595,fifo_intf_595,cstatus_csv_dumper_595);
    fifo_csv_dumper_596 = new("./depth596.csv");
    cstatus_csv_dumper_596 = new("./chan_status596.csv");
    fifo_monitor_596 = new(fifo_csv_dumper_596,fifo_intf_596,cstatus_csv_dumper_596);
    fifo_csv_dumper_597 = new("./depth597.csv");
    cstatus_csv_dumper_597 = new("./chan_status597.csv");
    fifo_monitor_597 = new(fifo_csv_dumper_597,fifo_intf_597,cstatus_csv_dumper_597);
    fifo_csv_dumper_598 = new("./depth598.csv");
    cstatus_csv_dumper_598 = new("./chan_status598.csv");
    fifo_monitor_598 = new(fifo_csv_dumper_598,fifo_intf_598,cstatus_csv_dumper_598);
    fifo_csv_dumper_599 = new("./depth599.csv");
    cstatus_csv_dumper_599 = new("./chan_status599.csv");
    fifo_monitor_599 = new(fifo_csv_dumper_599,fifo_intf_599,cstatus_csv_dumper_599);
    fifo_csv_dumper_600 = new("./depth600.csv");
    cstatus_csv_dumper_600 = new("./chan_status600.csv");
    fifo_monitor_600 = new(fifo_csv_dumper_600,fifo_intf_600,cstatus_csv_dumper_600);
    fifo_csv_dumper_601 = new("./depth601.csv");
    cstatus_csv_dumper_601 = new("./chan_status601.csv");
    fifo_monitor_601 = new(fifo_csv_dumper_601,fifo_intf_601,cstatus_csv_dumper_601);
    fifo_csv_dumper_602 = new("./depth602.csv");
    cstatus_csv_dumper_602 = new("./chan_status602.csv");
    fifo_monitor_602 = new(fifo_csv_dumper_602,fifo_intf_602,cstatus_csv_dumper_602);
    fifo_csv_dumper_603 = new("./depth603.csv");
    cstatus_csv_dumper_603 = new("./chan_status603.csv");
    fifo_monitor_603 = new(fifo_csv_dumper_603,fifo_intf_603,cstatus_csv_dumper_603);
    fifo_csv_dumper_604 = new("./depth604.csv");
    cstatus_csv_dumper_604 = new("./chan_status604.csv");
    fifo_monitor_604 = new(fifo_csv_dumper_604,fifo_intf_604,cstatus_csv_dumper_604);
    fifo_csv_dumper_605 = new("./depth605.csv");
    cstatus_csv_dumper_605 = new("./chan_status605.csv");
    fifo_monitor_605 = new(fifo_csv_dumper_605,fifo_intf_605,cstatus_csv_dumper_605);
    fifo_csv_dumper_606 = new("./depth606.csv");
    cstatus_csv_dumper_606 = new("./chan_status606.csv");
    fifo_monitor_606 = new(fifo_csv_dumper_606,fifo_intf_606,cstatus_csv_dumper_606);
    fifo_csv_dumper_607 = new("./depth607.csv");
    cstatus_csv_dumper_607 = new("./chan_status607.csv");
    fifo_monitor_607 = new(fifo_csv_dumper_607,fifo_intf_607,cstatus_csv_dumper_607);
    fifo_csv_dumper_608 = new("./depth608.csv");
    cstatus_csv_dumper_608 = new("./chan_status608.csv");
    fifo_monitor_608 = new(fifo_csv_dumper_608,fifo_intf_608,cstatus_csv_dumper_608);
    fifo_csv_dumper_609 = new("./depth609.csv");
    cstatus_csv_dumper_609 = new("./chan_status609.csv");
    fifo_monitor_609 = new(fifo_csv_dumper_609,fifo_intf_609,cstatus_csv_dumper_609);
    fifo_csv_dumper_610 = new("./depth610.csv");
    cstatus_csv_dumper_610 = new("./chan_status610.csv");
    fifo_monitor_610 = new(fifo_csv_dumper_610,fifo_intf_610,cstatus_csv_dumper_610);
    fifo_csv_dumper_611 = new("./depth611.csv");
    cstatus_csv_dumper_611 = new("./chan_status611.csv");
    fifo_monitor_611 = new(fifo_csv_dumper_611,fifo_intf_611,cstatus_csv_dumper_611);
    fifo_csv_dumper_612 = new("./depth612.csv");
    cstatus_csv_dumper_612 = new("./chan_status612.csv");
    fifo_monitor_612 = new(fifo_csv_dumper_612,fifo_intf_612,cstatus_csv_dumper_612);
    fifo_csv_dumper_613 = new("./depth613.csv");
    cstatus_csv_dumper_613 = new("./chan_status613.csv");
    fifo_monitor_613 = new(fifo_csv_dumper_613,fifo_intf_613,cstatus_csv_dumper_613);
    fifo_csv_dumper_614 = new("./depth614.csv");
    cstatus_csv_dumper_614 = new("./chan_status614.csv");
    fifo_monitor_614 = new(fifo_csv_dumper_614,fifo_intf_614,cstatus_csv_dumper_614);
    fifo_csv_dumper_615 = new("./depth615.csv");
    cstatus_csv_dumper_615 = new("./chan_status615.csv");
    fifo_monitor_615 = new(fifo_csv_dumper_615,fifo_intf_615,cstatus_csv_dumper_615);
    fifo_csv_dumper_616 = new("./depth616.csv");
    cstatus_csv_dumper_616 = new("./chan_status616.csv");
    fifo_monitor_616 = new(fifo_csv_dumper_616,fifo_intf_616,cstatus_csv_dumper_616);
    fifo_csv_dumper_617 = new("./depth617.csv");
    cstatus_csv_dumper_617 = new("./chan_status617.csv");
    fifo_monitor_617 = new(fifo_csv_dumper_617,fifo_intf_617,cstatus_csv_dumper_617);
    fifo_csv_dumper_618 = new("./depth618.csv");
    cstatus_csv_dumper_618 = new("./chan_status618.csv");
    fifo_monitor_618 = new(fifo_csv_dumper_618,fifo_intf_618,cstatus_csv_dumper_618);
    fifo_csv_dumper_619 = new("./depth619.csv");
    cstatus_csv_dumper_619 = new("./chan_status619.csv");
    fifo_monitor_619 = new(fifo_csv_dumper_619,fifo_intf_619,cstatus_csv_dumper_619);
    fifo_csv_dumper_620 = new("./depth620.csv");
    cstatus_csv_dumper_620 = new("./chan_status620.csv");
    fifo_monitor_620 = new(fifo_csv_dumper_620,fifo_intf_620,cstatus_csv_dumper_620);
    fifo_csv_dumper_621 = new("./depth621.csv");
    cstatus_csv_dumper_621 = new("./chan_status621.csv");
    fifo_monitor_621 = new(fifo_csv_dumper_621,fifo_intf_621,cstatus_csv_dumper_621);
    fifo_csv_dumper_622 = new("./depth622.csv");
    cstatus_csv_dumper_622 = new("./chan_status622.csv");
    fifo_monitor_622 = new(fifo_csv_dumper_622,fifo_intf_622,cstatus_csv_dumper_622);
    fifo_csv_dumper_623 = new("./depth623.csv");
    cstatus_csv_dumper_623 = new("./chan_status623.csv");
    fifo_monitor_623 = new(fifo_csv_dumper_623,fifo_intf_623,cstatus_csv_dumper_623);
    fifo_csv_dumper_624 = new("./depth624.csv");
    cstatus_csv_dumper_624 = new("./chan_status624.csv");
    fifo_monitor_624 = new(fifo_csv_dumper_624,fifo_intf_624,cstatus_csv_dumper_624);
    fifo_csv_dumper_625 = new("./depth625.csv");
    cstatus_csv_dumper_625 = new("./chan_status625.csv");
    fifo_monitor_625 = new(fifo_csv_dumper_625,fifo_intf_625,cstatus_csv_dumper_625);
    fifo_csv_dumper_626 = new("./depth626.csv");
    cstatus_csv_dumper_626 = new("./chan_status626.csv");
    fifo_monitor_626 = new(fifo_csv_dumper_626,fifo_intf_626,cstatus_csv_dumper_626);
    fifo_csv_dumper_627 = new("./depth627.csv");
    cstatus_csv_dumper_627 = new("./chan_status627.csv");
    fifo_monitor_627 = new(fifo_csv_dumper_627,fifo_intf_627,cstatus_csv_dumper_627);
    fifo_csv_dumper_628 = new("./depth628.csv");
    cstatus_csv_dumper_628 = new("./chan_status628.csv");
    fifo_monitor_628 = new(fifo_csv_dumper_628,fifo_intf_628,cstatus_csv_dumper_628);
    fifo_csv_dumper_629 = new("./depth629.csv");
    cstatus_csv_dumper_629 = new("./chan_status629.csv");
    fifo_monitor_629 = new(fifo_csv_dumper_629,fifo_intf_629,cstatus_csv_dumper_629);
    fifo_csv_dumper_630 = new("./depth630.csv");
    cstatus_csv_dumper_630 = new("./chan_status630.csv");
    fifo_monitor_630 = new(fifo_csv_dumper_630,fifo_intf_630,cstatus_csv_dumper_630);
    fifo_csv_dumper_631 = new("./depth631.csv");
    cstatus_csv_dumper_631 = new("./chan_status631.csv");
    fifo_monitor_631 = new(fifo_csv_dumper_631,fifo_intf_631,cstatus_csv_dumper_631);
    fifo_csv_dumper_632 = new("./depth632.csv");
    cstatus_csv_dumper_632 = new("./chan_status632.csv");
    fifo_monitor_632 = new(fifo_csv_dumper_632,fifo_intf_632,cstatus_csv_dumper_632);
    fifo_csv_dumper_633 = new("./depth633.csv");
    cstatus_csv_dumper_633 = new("./chan_status633.csv");
    fifo_monitor_633 = new(fifo_csv_dumper_633,fifo_intf_633,cstatus_csv_dumper_633);
    fifo_csv_dumper_634 = new("./depth634.csv");
    cstatus_csv_dumper_634 = new("./chan_status634.csv");
    fifo_monitor_634 = new(fifo_csv_dumper_634,fifo_intf_634,cstatus_csv_dumper_634);
    fifo_csv_dumper_635 = new("./depth635.csv");
    cstatus_csv_dumper_635 = new("./chan_status635.csv");
    fifo_monitor_635 = new(fifo_csv_dumper_635,fifo_intf_635,cstatus_csv_dumper_635);
    fifo_csv_dumper_636 = new("./depth636.csv");
    cstatus_csv_dumper_636 = new("./chan_status636.csv");
    fifo_monitor_636 = new(fifo_csv_dumper_636,fifo_intf_636,cstatus_csv_dumper_636);
    fifo_csv_dumper_637 = new("./depth637.csv");
    cstatus_csv_dumper_637 = new("./chan_status637.csv");
    fifo_monitor_637 = new(fifo_csv_dumper_637,fifo_intf_637,cstatus_csv_dumper_637);
    fifo_csv_dumper_638 = new("./depth638.csv");
    cstatus_csv_dumper_638 = new("./chan_status638.csv");
    fifo_monitor_638 = new(fifo_csv_dumper_638,fifo_intf_638,cstatus_csv_dumper_638);
    fifo_csv_dumper_639 = new("./depth639.csv");
    cstatus_csv_dumper_639 = new("./chan_status639.csv");
    fifo_monitor_639 = new(fifo_csv_dumper_639,fifo_intf_639,cstatus_csv_dumper_639);
    fifo_csv_dumper_640 = new("./depth640.csv");
    cstatus_csv_dumper_640 = new("./chan_status640.csv");
    fifo_monitor_640 = new(fifo_csv_dumper_640,fifo_intf_640,cstatus_csv_dumper_640);
    fifo_csv_dumper_641 = new("./depth641.csv");
    cstatus_csv_dumper_641 = new("./chan_status641.csv");
    fifo_monitor_641 = new(fifo_csv_dumper_641,fifo_intf_641,cstatus_csv_dumper_641);
    fifo_csv_dumper_642 = new("./depth642.csv");
    cstatus_csv_dumper_642 = new("./chan_status642.csv");
    fifo_monitor_642 = new(fifo_csv_dumper_642,fifo_intf_642,cstatus_csv_dumper_642);
    fifo_csv_dumper_643 = new("./depth643.csv");
    cstatus_csv_dumper_643 = new("./chan_status643.csv");
    fifo_monitor_643 = new(fifo_csv_dumper_643,fifo_intf_643,cstatus_csv_dumper_643);
    fifo_csv_dumper_644 = new("./depth644.csv");
    cstatus_csv_dumper_644 = new("./chan_status644.csv");
    fifo_monitor_644 = new(fifo_csv_dumper_644,fifo_intf_644,cstatus_csv_dumper_644);
    fifo_csv_dumper_645 = new("./depth645.csv");
    cstatus_csv_dumper_645 = new("./chan_status645.csv");
    fifo_monitor_645 = new(fifo_csv_dumper_645,fifo_intf_645,cstatus_csv_dumper_645);
    fifo_csv_dumper_646 = new("./depth646.csv");
    cstatus_csv_dumper_646 = new("./chan_status646.csv");
    fifo_monitor_646 = new(fifo_csv_dumper_646,fifo_intf_646,cstatus_csv_dumper_646);
    fifo_csv_dumper_647 = new("./depth647.csv");
    cstatus_csv_dumper_647 = new("./chan_status647.csv");
    fifo_monitor_647 = new(fifo_csv_dumper_647,fifo_intf_647,cstatus_csv_dumper_647);
    fifo_csv_dumper_648 = new("./depth648.csv");
    cstatus_csv_dumper_648 = new("./chan_status648.csv");
    fifo_monitor_648 = new(fifo_csv_dumper_648,fifo_intf_648,cstatus_csv_dumper_648);
    fifo_csv_dumper_649 = new("./depth649.csv");
    cstatus_csv_dumper_649 = new("./chan_status649.csv");
    fifo_monitor_649 = new(fifo_csv_dumper_649,fifo_intf_649,cstatus_csv_dumper_649);
    fifo_csv_dumper_650 = new("./depth650.csv");
    cstatus_csv_dumper_650 = new("./chan_status650.csv");
    fifo_monitor_650 = new(fifo_csv_dumper_650,fifo_intf_650,cstatus_csv_dumper_650);
    fifo_csv_dumper_651 = new("./depth651.csv");
    cstatus_csv_dumper_651 = new("./chan_status651.csv");
    fifo_monitor_651 = new(fifo_csv_dumper_651,fifo_intf_651,cstatus_csv_dumper_651);
    fifo_csv_dumper_652 = new("./depth652.csv");
    cstatus_csv_dumper_652 = new("./chan_status652.csv");
    fifo_monitor_652 = new(fifo_csv_dumper_652,fifo_intf_652,cstatus_csv_dumper_652);
    fifo_csv_dumper_653 = new("./depth653.csv");
    cstatus_csv_dumper_653 = new("./chan_status653.csv");
    fifo_monitor_653 = new(fifo_csv_dumper_653,fifo_intf_653,cstatus_csv_dumper_653);
    fifo_csv_dumper_654 = new("./depth654.csv");
    cstatus_csv_dumper_654 = new("./chan_status654.csv");
    fifo_monitor_654 = new(fifo_csv_dumper_654,fifo_intf_654,cstatus_csv_dumper_654);
    fifo_csv_dumper_655 = new("./depth655.csv");
    cstatus_csv_dumper_655 = new("./chan_status655.csv");
    fifo_monitor_655 = new(fifo_csv_dumper_655,fifo_intf_655,cstatus_csv_dumper_655);
    fifo_csv_dumper_656 = new("./depth656.csv");
    cstatus_csv_dumper_656 = new("./chan_status656.csv");
    fifo_monitor_656 = new(fifo_csv_dumper_656,fifo_intf_656,cstatus_csv_dumper_656);
    fifo_csv_dumper_657 = new("./depth657.csv");
    cstatus_csv_dumper_657 = new("./chan_status657.csv");
    fifo_monitor_657 = new(fifo_csv_dumper_657,fifo_intf_657,cstatus_csv_dumper_657);
    fifo_csv_dumper_658 = new("./depth658.csv");
    cstatus_csv_dumper_658 = new("./chan_status658.csv");
    fifo_monitor_658 = new(fifo_csv_dumper_658,fifo_intf_658,cstatus_csv_dumper_658);
    fifo_csv_dumper_659 = new("./depth659.csv");
    cstatus_csv_dumper_659 = new("./chan_status659.csv");
    fifo_monitor_659 = new(fifo_csv_dumper_659,fifo_intf_659,cstatus_csv_dumper_659);
    fifo_csv_dumper_660 = new("./depth660.csv");
    cstatus_csv_dumper_660 = new("./chan_status660.csv");
    fifo_monitor_660 = new(fifo_csv_dumper_660,fifo_intf_660,cstatus_csv_dumper_660);
    fifo_csv_dumper_661 = new("./depth661.csv");
    cstatus_csv_dumper_661 = new("./chan_status661.csv");
    fifo_monitor_661 = new(fifo_csv_dumper_661,fifo_intf_661,cstatus_csv_dumper_661);
    fifo_csv_dumper_662 = new("./depth662.csv");
    cstatus_csv_dumper_662 = new("./chan_status662.csv");
    fifo_monitor_662 = new(fifo_csv_dumper_662,fifo_intf_662,cstatus_csv_dumper_662);
    fifo_csv_dumper_663 = new("./depth663.csv");
    cstatus_csv_dumper_663 = new("./chan_status663.csv");
    fifo_monitor_663 = new(fifo_csv_dumper_663,fifo_intf_663,cstatus_csv_dumper_663);
    fifo_csv_dumper_664 = new("./depth664.csv");
    cstatus_csv_dumper_664 = new("./chan_status664.csv");
    fifo_monitor_664 = new(fifo_csv_dumper_664,fifo_intf_664,cstatus_csv_dumper_664);
    fifo_csv_dumper_665 = new("./depth665.csv");
    cstatus_csv_dumper_665 = new("./chan_status665.csv");
    fifo_monitor_665 = new(fifo_csv_dumper_665,fifo_intf_665,cstatus_csv_dumper_665);
    fifo_csv_dumper_666 = new("./depth666.csv");
    cstatus_csv_dumper_666 = new("./chan_status666.csv");
    fifo_monitor_666 = new(fifo_csv_dumper_666,fifo_intf_666,cstatus_csv_dumper_666);
    fifo_csv_dumper_667 = new("./depth667.csv");
    cstatus_csv_dumper_667 = new("./chan_status667.csv");
    fifo_monitor_667 = new(fifo_csv_dumper_667,fifo_intf_667,cstatus_csv_dumper_667);
    fifo_csv_dumper_668 = new("./depth668.csv");
    cstatus_csv_dumper_668 = new("./chan_status668.csv");
    fifo_monitor_668 = new(fifo_csv_dumper_668,fifo_intf_668,cstatus_csv_dumper_668);
    fifo_csv_dumper_669 = new("./depth669.csv");
    cstatus_csv_dumper_669 = new("./chan_status669.csv");
    fifo_monitor_669 = new(fifo_csv_dumper_669,fifo_intf_669,cstatus_csv_dumper_669);
    fifo_csv_dumper_670 = new("./depth670.csv");
    cstatus_csv_dumper_670 = new("./chan_status670.csv");
    fifo_monitor_670 = new(fifo_csv_dumper_670,fifo_intf_670,cstatus_csv_dumper_670);
    fifo_csv_dumper_671 = new("./depth671.csv");
    cstatus_csv_dumper_671 = new("./chan_status671.csv");
    fifo_monitor_671 = new(fifo_csv_dumper_671,fifo_intf_671,cstatus_csv_dumper_671);
    fifo_csv_dumper_672 = new("./depth672.csv");
    cstatus_csv_dumper_672 = new("./chan_status672.csv");
    fifo_monitor_672 = new(fifo_csv_dumper_672,fifo_intf_672,cstatus_csv_dumper_672);
    fifo_csv_dumper_673 = new("./depth673.csv");
    cstatus_csv_dumper_673 = new("./chan_status673.csv");
    fifo_monitor_673 = new(fifo_csv_dumper_673,fifo_intf_673,cstatus_csv_dumper_673);
    fifo_csv_dumper_674 = new("./depth674.csv");
    cstatus_csv_dumper_674 = new("./chan_status674.csv");
    fifo_monitor_674 = new(fifo_csv_dumper_674,fifo_intf_674,cstatus_csv_dumper_674);
    fifo_csv_dumper_675 = new("./depth675.csv");
    cstatus_csv_dumper_675 = new("./chan_status675.csv");
    fifo_monitor_675 = new(fifo_csv_dumper_675,fifo_intf_675,cstatus_csv_dumper_675);
    fifo_csv_dumper_676 = new("./depth676.csv");
    cstatus_csv_dumper_676 = new("./chan_status676.csv");
    fifo_monitor_676 = new(fifo_csv_dumper_676,fifo_intf_676,cstatus_csv_dumper_676);
    fifo_csv_dumper_677 = new("./depth677.csv");
    cstatus_csv_dumper_677 = new("./chan_status677.csv");
    fifo_monitor_677 = new(fifo_csv_dumper_677,fifo_intf_677,cstatus_csv_dumper_677);
    fifo_csv_dumper_678 = new("./depth678.csv");
    cstatus_csv_dumper_678 = new("./chan_status678.csv");
    fifo_monitor_678 = new(fifo_csv_dumper_678,fifo_intf_678,cstatus_csv_dumper_678);
    fifo_csv_dumper_679 = new("./depth679.csv");
    cstatus_csv_dumper_679 = new("./chan_status679.csv");
    fifo_monitor_679 = new(fifo_csv_dumper_679,fifo_intf_679,cstatus_csv_dumper_679);
    fifo_csv_dumper_680 = new("./depth680.csv");
    cstatus_csv_dumper_680 = new("./chan_status680.csv");
    fifo_monitor_680 = new(fifo_csv_dumper_680,fifo_intf_680,cstatus_csv_dumper_680);
    fifo_csv_dumper_681 = new("./depth681.csv");
    cstatus_csv_dumper_681 = new("./chan_status681.csv");
    fifo_monitor_681 = new(fifo_csv_dumper_681,fifo_intf_681,cstatus_csv_dumper_681);
    fifo_csv_dumper_682 = new("./depth682.csv");
    cstatus_csv_dumper_682 = new("./chan_status682.csv");
    fifo_monitor_682 = new(fifo_csv_dumper_682,fifo_intf_682,cstatus_csv_dumper_682);
    fifo_csv_dumper_683 = new("./depth683.csv");
    cstatus_csv_dumper_683 = new("./chan_status683.csv");
    fifo_monitor_683 = new(fifo_csv_dumper_683,fifo_intf_683,cstatus_csv_dumper_683);
    fifo_csv_dumper_684 = new("./depth684.csv");
    cstatus_csv_dumper_684 = new("./chan_status684.csv");
    fifo_monitor_684 = new(fifo_csv_dumper_684,fifo_intf_684,cstatus_csv_dumper_684);
    fifo_csv_dumper_685 = new("./depth685.csv");
    cstatus_csv_dumper_685 = new("./chan_status685.csv");
    fifo_monitor_685 = new(fifo_csv_dumper_685,fifo_intf_685,cstatus_csv_dumper_685);
    fifo_csv_dumper_686 = new("./depth686.csv");
    cstatus_csv_dumper_686 = new("./chan_status686.csv");
    fifo_monitor_686 = new(fifo_csv_dumper_686,fifo_intf_686,cstatus_csv_dumper_686);
    fifo_csv_dumper_687 = new("./depth687.csv");
    cstatus_csv_dumper_687 = new("./chan_status687.csv");
    fifo_monitor_687 = new(fifo_csv_dumper_687,fifo_intf_687,cstatus_csv_dumper_687);
    fifo_csv_dumper_688 = new("./depth688.csv");
    cstatus_csv_dumper_688 = new("./chan_status688.csv");
    fifo_monitor_688 = new(fifo_csv_dumper_688,fifo_intf_688,cstatus_csv_dumper_688);
    fifo_csv_dumper_689 = new("./depth689.csv");
    cstatus_csv_dumper_689 = new("./chan_status689.csv");
    fifo_monitor_689 = new(fifo_csv_dumper_689,fifo_intf_689,cstatus_csv_dumper_689);
    fifo_csv_dumper_690 = new("./depth690.csv");
    cstatus_csv_dumper_690 = new("./chan_status690.csv");
    fifo_monitor_690 = new(fifo_csv_dumper_690,fifo_intf_690,cstatus_csv_dumper_690);
    fifo_csv_dumper_691 = new("./depth691.csv");
    cstatus_csv_dumper_691 = new("./chan_status691.csv");
    fifo_monitor_691 = new(fifo_csv_dumper_691,fifo_intf_691,cstatus_csv_dumper_691);
    fifo_csv_dumper_692 = new("./depth692.csv");
    cstatus_csv_dumper_692 = new("./chan_status692.csv");
    fifo_monitor_692 = new(fifo_csv_dumper_692,fifo_intf_692,cstatus_csv_dumper_692);
    fifo_csv_dumper_693 = new("./depth693.csv");
    cstatus_csv_dumper_693 = new("./chan_status693.csv");
    fifo_monitor_693 = new(fifo_csv_dumper_693,fifo_intf_693,cstatus_csv_dumper_693);
    fifo_csv_dumper_694 = new("./depth694.csv");
    cstatus_csv_dumper_694 = new("./chan_status694.csv");
    fifo_monitor_694 = new(fifo_csv_dumper_694,fifo_intf_694,cstatus_csv_dumper_694);
    fifo_csv_dumper_695 = new("./depth695.csv");
    cstatus_csv_dumper_695 = new("./chan_status695.csv");
    fifo_monitor_695 = new(fifo_csv_dumper_695,fifo_intf_695,cstatus_csv_dumper_695);
    fifo_csv_dumper_696 = new("./depth696.csv");
    cstatus_csv_dumper_696 = new("./chan_status696.csv");
    fifo_monitor_696 = new(fifo_csv_dumper_696,fifo_intf_696,cstatus_csv_dumper_696);
    fifo_csv_dumper_697 = new("./depth697.csv");
    cstatus_csv_dumper_697 = new("./chan_status697.csv");
    fifo_monitor_697 = new(fifo_csv_dumper_697,fifo_intf_697,cstatus_csv_dumper_697);
    fifo_csv_dumper_698 = new("./depth698.csv");
    cstatus_csv_dumper_698 = new("./chan_status698.csv");
    fifo_monitor_698 = new(fifo_csv_dumper_698,fifo_intf_698,cstatus_csv_dumper_698);
    fifo_csv_dumper_699 = new("./depth699.csv");
    cstatus_csv_dumper_699 = new("./chan_status699.csv");
    fifo_monitor_699 = new(fifo_csv_dumper_699,fifo_intf_699,cstatus_csv_dumper_699);
    fifo_csv_dumper_700 = new("./depth700.csv");
    cstatus_csv_dumper_700 = new("./chan_status700.csv");
    fifo_monitor_700 = new(fifo_csv_dumper_700,fifo_intf_700,cstatus_csv_dumper_700);
    fifo_csv_dumper_701 = new("./depth701.csv");
    cstatus_csv_dumper_701 = new("./chan_status701.csv");
    fifo_monitor_701 = new(fifo_csv_dumper_701,fifo_intf_701,cstatus_csv_dumper_701);
    fifo_csv_dumper_702 = new("./depth702.csv");
    cstatus_csv_dumper_702 = new("./chan_status702.csv");
    fifo_monitor_702 = new(fifo_csv_dumper_702,fifo_intf_702,cstatus_csv_dumper_702);
    fifo_csv_dumper_703 = new("./depth703.csv");
    cstatus_csv_dumper_703 = new("./chan_status703.csv");
    fifo_monitor_703 = new(fifo_csv_dumper_703,fifo_intf_703,cstatus_csv_dumper_703);
    fifo_csv_dumper_704 = new("./depth704.csv");
    cstatus_csv_dumper_704 = new("./chan_status704.csv");
    fifo_monitor_704 = new(fifo_csv_dumper_704,fifo_intf_704,cstatus_csv_dumper_704);
    fifo_csv_dumper_705 = new("./depth705.csv");
    cstatus_csv_dumper_705 = new("./chan_status705.csv");
    fifo_monitor_705 = new(fifo_csv_dumper_705,fifo_intf_705,cstatus_csv_dumper_705);
    fifo_csv_dumper_706 = new("./depth706.csv");
    cstatus_csv_dumper_706 = new("./chan_status706.csv");
    fifo_monitor_706 = new(fifo_csv_dumper_706,fifo_intf_706,cstatus_csv_dumper_706);
    fifo_csv_dumper_707 = new("./depth707.csv");
    cstatus_csv_dumper_707 = new("./chan_status707.csv");
    fifo_monitor_707 = new(fifo_csv_dumper_707,fifo_intf_707,cstatus_csv_dumper_707);
    fifo_csv_dumper_708 = new("./depth708.csv");
    cstatus_csv_dumper_708 = new("./chan_status708.csv");
    fifo_monitor_708 = new(fifo_csv_dumper_708,fifo_intf_708,cstatus_csv_dumper_708);
    fifo_csv_dumper_709 = new("./depth709.csv");
    cstatus_csv_dumper_709 = new("./chan_status709.csv");
    fifo_monitor_709 = new(fifo_csv_dumper_709,fifo_intf_709,cstatus_csv_dumper_709);
    fifo_csv_dumper_710 = new("./depth710.csv");
    cstatus_csv_dumper_710 = new("./chan_status710.csv");
    fifo_monitor_710 = new(fifo_csv_dumper_710,fifo_intf_710,cstatus_csv_dumper_710);
    fifo_csv_dumper_711 = new("./depth711.csv");
    cstatus_csv_dumper_711 = new("./chan_status711.csv");
    fifo_monitor_711 = new(fifo_csv_dumper_711,fifo_intf_711,cstatus_csv_dumper_711);
    fifo_csv_dumper_712 = new("./depth712.csv");
    cstatus_csv_dumper_712 = new("./chan_status712.csv");
    fifo_monitor_712 = new(fifo_csv_dumper_712,fifo_intf_712,cstatus_csv_dumper_712);
    fifo_csv_dumper_713 = new("./depth713.csv");
    cstatus_csv_dumper_713 = new("./chan_status713.csv");
    fifo_monitor_713 = new(fifo_csv_dumper_713,fifo_intf_713,cstatus_csv_dumper_713);
    fifo_csv_dumper_714 = new("./depth714.csv");
    cstatus_csv_dumper_714 = new("./chan_status714.csv");
    fifo_monitor_714 = new(fifo_csv_dumper_714,fifo_intf_714,cstatus_csv_dumper_714);
    fifo_csv_dumper_715 = new("./depth715.csv");
    cstatus_csv_dumper_715 = new("./chan_status715.csv");
    fifo_monitor_715 = new(fifo_csv_dumper_715,fifo_intf_715,cstatus_csv_dumper_715);
    fifo_csv_dumper_716 = new("./depth716.csv");
    cstatus_csv_dumper_716 = new("./chan_status716.csv");
    fifo_monitor_716 = new(fifo_csv_dumper_716,fifo_intf_716,cstatus_csv_dumper_716);
    fifo_csv_dumper_717 = new("./depth717.csv");
    cstatus_csv_dumper_717 = new("./chan_status717.csv");
    fifo_monitor_717 = new(fifo_csv_dumper_717,fifo_intf_717,cstatus_csv_dumper_717);
    fifo_csv_dumper_718 = new("./depth718.csv");
    cstatus_csv_dumper_718 = new("./chan_status718.csv");
    fifo_monitor_718 = new(fifo_csv_dumper_718,fifo_intf_718,cstatus_csv_dumper_718);
    fifo_csv_dumper_719 = new("./depth719.csv");
    cstatus_csv_dumper_719 = new("./chan_status719.csv");
    fifo_monitor_719 = new(fifo_csv_dumper_719,fifo_intf_719,cstatus_csv_dumper_719);
    fifo_csv_dumper_720 = new("./depth720.csv");
    cstatus_csv_dumper_720 = new("./chan_status720.csv");
    fifo_monitor_720 = new(fifo_csv_dumper_720,fifo_intf_720,cstatus_csv_dumper_720);
    fifo_csv_dumper_721 = new("./depth721.csv");
    cstatus_csv_dumper_721 = new("./chan_status721.csv");
    fifo_monitor_721 = new(fifo_csv_dumper_721,fifo_intf_721,cstatus_csv_dumper_721);
    fifo_csv_dumper_722 = new("./depth722.csv");
    cstatus_csv_dumper_722 = new("./chan_status722.csv");
    fifo_monitor_722 = new(fifo_csv_dumper_722,fifo_intf_722,cstatus_csv_dumper_722);
    fifo_csv_dumper_723 = new("./depth723.csv");
    cstatus_csv_dumper_723 = new("./chan_status723.csv");
    fifo_monitor_723 = new(fifo_csv_dumper_723,fifo_intf_723,cstatus_csv_dumper_723);
    fifo_csv_dumper_724 = new("./depth724.csv");
    cstatus_csv_dumper_724 = new("./chan_status724.csv");
    fifo_monitor_724 = new(fifo_csv_dumper_724,fifo_intf_724,cstatus_csv_dumper_724);
    fifo_csv_dumper_725 = new("./depth725.csv");
    cstatus_csv_dumper_725 = new("./chan_status725.csv");
    fifo_monitor_725 = new(fifo_csv_dumper_725,fifo_intf_725,cstatus_csv_dumper_725);
    fifo_csv_dumper_726 = new("./depth726.csv");
    cstatus_csv_dumper_726 = new("./chan_status726.csv");
    fifo_monitor_726 = new(fifo_csv_dumper_726,fifo_intf_726,cstatus_csv_dumper_726);
    fifo_csv_dumper_727 = new("./depth727.csv");
    cstatus_csv_dumper_727 = new("./chan_status727.csv");
    fifo_monitor_727 = new(fifo_csv_dumper_727,fifo_intf_727,cstatus_csv_dumper_727);
    fifo_csv_dumper_728 = new("./depth728.csv");
    cstatus_csv_dumper_728 = new("./chan_status728.csv");
    fifo_monitor_728 = new(fifo_csv_dumper_728,fifo_intf_728,cstatus_csv_dumper_728);
    fifo_csv_dumper_729 = new("./depth729.csv");
    cstatus_csv_dumper_729 = new("./chan_status729.csv");
    fifo_monitor_729 = new(fifo_csv_dumper_729,fifo_intf_729,cstatus_csv_dumper_729);
    fifo_csv_dumper_730 = new("./depth730.csv");
    cstatus_csv_dumper_730 = new("./chan_status730.csv");
    fifo_monitor_730 = new(fifo_csv_dumper_730,fifo_intf_730,cstatus_csv_dumper_730);
    fifo_csv_dumper_731 = new("./depth731.csv");
    cstatus_csv_dumper_731 = new("./chan_status731.csv");
    fifo_monitor_731 = new(fifo_csv_dumper_731,fifo_intf_731,cstatus_csv_dumper_731);
    fifo_csv_dumper_732 = new("./depth732.csv");
    cstatus_csv_dumper_732 = new("./chan_status732.csv");
    fifo_monitor_732 = new(fifo_csv_dumper_732,fifo_intf_732,cstatus_csv_dumper_732);
    fifo_csv_dumper_733 = new("./depth733.csv");
    cstatus_csv_dumper_733 = new("./chan_status733.csv");
    fifo_monitor_733 = new(fifo_csv_dumper_733,fifo_intf_733,cstatus_csv_dumper_733);
    fifo_csv_dumper_734 = new("./depth734.csv");
    cstatus_csv_dumper_734 = new("./chan_status734.csv");
    fifo_monitor_734 = new(fifo_csv_dumper_734,fifo_intf_734,cstatus_csv_dumper_734);
    fifo_csv_dumper_735 = new("./depth735.csv");
    cstatus_csv_dumper_735 = new("./chan_status735.csv");
    fifo_monitor_735 = new(fifo_csv_dumper_735,fifo_intf_735,cstatus_csv_dumper_735);
    fifo_csv_dumper_736 = new("./depth736.csv");
    cstatus_csv_dumper_736 = new("./chan_status736.csv");
    fifo_monitor_736 = new(fifo_csv_dumper_736,fifo_intf_736,cstatus_csv_dumper_736);
    fifo_csv_dumper_737 = new("./depth737.csv");
    cstatus_csv_dumper_737 = new("./chan_status737.csv");
    fifo_monitor_737 = new(fifo_csv_dumper_737,fifo_intf_737,cstatus_csv_dumper_737);
    fifo_csv_dumper_738 = new("./depth738.csv");
    cstatus_csv_dumper_738 = new("./chan_status738.csv");
    fifo_monitor_738 = new(fifo_csv_dumper_738,fifo_intf_738,cstatus_csv_dumper_738);
    fifo_csv_dumper_739 = new("./depth739.csv");
    cstatus_csv_dumper_739 = new("./chan_status739.csv");
    fifo_monitor_739 = new(fifo_csv_dumper_739,fifo_intf_739,cstatus_csv_dumper_739);
    fifo_csv_dumper_740 = new("./depth740.csv");
    cstatus_csv_dumper_740 = new("./chan_status740.csv");
    fifo_monitor_740 = new(fifo_csv_dumper_740,fifo_intf_740,cstatus_csv_dumper_740);
    fifo_csv_dumper_741 = new("./depth741.csv");
    cstatus_csv_dumper_741 = new("./chan_status741.csv");
    fifo_monitor_741 = new(fifo_csv_dumper_741,fifo_intf_741,cstatus_csv_dumper_741);
    fifo_csv_dumper_742 = new("./depth742.csv");
    cstatus_csv_dumper_742 = new("./chan_status742.csv");
    fifo_monitor_742 = new(fifo_csv_dumper_742,fifo_intf_742,cstatus_csv_dumper_742);
    fifo_csv_dumper_743 = new("./depth743.csv");
    cstatus_csv_dumper_743 = new("./chan_status743.csv");
    fifo_monitor_743 = new(fifo_csv_dumper_743,fifo_intf_743,cstatus_csv_dumper_743);
    fifo_csv_dumper_744 = new("./depth744.csv");
    cstatus_csv_dumper_744 = new("./chan_status744.csv");
    fifo_monitor_744 = new(fifo_csv_dumper_744,fifo_intf_744,cstatus_csv_dumper_744);
    fifo_csv_dumper_745 = new("./depth745.csv");
    cstatus_csv_dumper_745 = new("./chan_status745.csv");
    fifo_monitor_745 = new(fifo_csv_dumper_745,fifo_intf_745,cstatus_csv_dumper_745);
    fifo_csv_dumper_746 = new("./depth746.csv");
    cstatus_csv_dumper_746 = new("./chan_status746.csv");
    fifo_monitor_746 = new(fifo_csv_dumper_746,fifo_intf_746,cstatus_csv_dumper_746);
    fifo_csv_dumper_747 = new("./depth747.csv");
    cstatus_csv_dumper_747 = new("./chan_status747.csv");
    fifo_monitor_747 = new(fifo_csv_dumper_747,fifo_intf_747,cstatus_csv_dumper_747);
    fifo_csv_dumper_748 = new("./depth748.csv");
    cstatus_csv_dumper_748 = new("./chan_status748.csv");
    fifo_monitor_748 = new(fifo_csv_dumper_748,fifo_intf_748,cstatus_csv_dumper_748);
    fifo_csv_dumper_749 = new("./depth749.csv");
    cstatus_csv_dumper_749 = new("./chan_status749.csv");
    fifo_monitor_749 = new(fifo_csv_dumper_749,fifo_intf_749,cstatus_csv_dumper_749);
    fifo_csv_dumper_750 = new("./depth750.csv");
    cstatus_csv_dumper_750 = new("./chan_status750.csv");
    fifo_monitor_750 = new(fifo_csv_dumper_750,fifo_intf_750,cstatus_csv_dumper_750);
    fifo_csv_dumper_751 = new("./depth751.csv");
    cstatus_csv_dumper_751 = new("./chan_status751.csv");
    fifo_monitor_751 = new(fifo_csv_dumper_751,fifo_intf_751,cstatus_csv_dumper_751);
    fifo_csv_dumper_752 = new("./depth752.csv");
    cstatus_csv_dumper_752 = new("./chan_status752.csv");
    fifo_monitor_752 = new(fifo_csv_dumper_752,fifo_intf_752,cstatus_csv_dumper_752);
    fifo_csv_dumper_753 = new("./depth753.csv");
    cstatus_csv_dumper_753 = new("./chan_status753.csv");
    fifo_monitor_753 = new(fifo_csv_dumper_753,fifo_intf_753,cstatus_csv_dumper_753);
    fifo_csv_dumper_754 = new("./depth754.csv");
    cstatus_csv_dumper_754 = new("./chan_status754.csv");
    fifo_monitor_754 = new(fifo_csv_dumper_754,fifo_intf_754,cstatus_csv_dumper_754);
    fifo_csv_dumper_755 = new("./depth755.csv");
    cstatus_csv_dumper_755 = new("./chan_status755.csv");
    fifo_monitor_755 = new(fifo_csv_dumper_755,fifo_intf_755,cstatus_csv_dumper_755);
    fifo_csv_dumper_756 = new("./depth756.csv");
    cstatus_csv_dumper_756 = new("./chan_status756.csv");
    fifo_monitor_756 = new(fifo_csv_dumper_756,fifo_intf_756,cstatus_csv_dumper_756);
    fifo_csv_dumper_757 = new("./depth757.csv");
    cstatus_csv_dumper_757 = new("./chan_status757.csv");
    fifo_monitor_757 = new(fifo_csv_dumper_757,fifo_intf_757,cstatus_csv_dumper_757);
    fifo_csv_dumper_758 = new("./depth758.csv");
    cstatus_csv_dumper_758 = new("./chan_status758.csv");
    fifo_monitor_758 = new(fifo_csv_dumper_758,fifo_intf_758,cstatus_csv_dumper_758);
    fifo_csv_dumper_759 = new("./depth759.csv");
    cstatus_csv_dumper_759 = new("./chan_status759.csv");
    fifo_monitor_759 = new(fifo_csv_dumper_759,fifo_intf_759,cstatus_csv_dumper_759);
    fifo_csv_dumper_760 = new("./depth760.csv");
    cstatus_csv_dumper_760 = new("./chan_status760.csv");
    fifo_monitor_760 = new(fifo_csv_dumper_760,fifo_intf_760,cstatus_csv_dumper_760);
    fifo_csv_dumper_761 = new("./depth761.csv");
    cstatus_csv_dumper_761 = new("./chan_status761.csv");
    fifo_monitor_761 = new(fifo_csv_dumper_761,fifo_intf_761,cstatus_csv_dumper_761);
    fifo_csv_dumper_762 = new("./depth762.csv");
    cstatus_csv_dumper_762 = new("./chan_status762.csv");
    fifo_monitor_762 = new(fifo_csv_dumper_762,fifo_intf_762,cstatus_csv_dumper_762);
    fifo_csv_dumper_763 = new("./depth763.csv");
    cstatus_csv_dumper_763 = new("./chan_status763.csv");
    fifo_monitor_763 = new(fifo_csv_dumper_763,fifo_intf_763,cstatus_csv_dumper_763);
    fifo_csv_dumper_764 = new("./depth764.csv");
    cstatus_csv_dumper_764 = new("./chan_status764.csv");
    fifo_monitor_764 = new(fifo_csv_dumper_764,fifo_intf_764,cstatus_csv_dumper_764);
    fifo_csv_dumper_765 = new("./depth765.csv");
    cstatus_csv_dumper_765 = new("./chan_status765.csv");
    fifo_monitor_765 = new(fifo_csv_dumper_765,fifo_intf_765,cstatus_csv_dumper_765);
    fifo_csv_dumper_766 = new("./depth766.csv");
    cstatus_csv_dumper_766 = new("./chan_status766.csv");
    fifo_monitor_766 = new(fifo_csv_dumper_766,fifo_intf_766,cstatus_csv_dumper_766);
    fifo_csv_dumper_767 = new("./depth767.csv");
    cstatus_csv_dumper_767 = new("./chan_status767.csv");
    fifo_monitor_767 = new(fifo_csv_dumper_767,fifo_intf_767,cstatus_csv_dumper_767);
    fifo_csv_dumper_768 = new("./depth768.csv");
    cstatus_csv_dumper_768 = new("./chan_status768.csv");
    fifo_monitor_768 = new(fifo_csv_dumper_768,fifo_intf_768,cstatus_csv_dumper_768);
    fifo_csv_dumper_769 = new("./depth769.csv");
    cstatus_csv_dumper_769 = new("./chan_status769.csv");
    fifo_monitor_769 = new(fifo_csv_dumper_769,fifo_intf_769,cstatus_csv_dumper_769);
    fifo_csv_dumper_770 = new("./depth770.csv");
    cstatus_csv_dumper_770 = new("./chan_status770.csv");
    fifo_monitor_770 = new(fifo_csv_dumper_770,fifo_intf_770,cstatus_csv_dumper_770);
    fifo_csv_dumper_771 = new("./depth771.csv");
    cstatus_csv_dumper_771 = new("./chan_status771.csv");
    fifo_monitor_771 = new(fifo_csv_dumper_771,fifo_intf_771,cstatus_csv_dumper_771);
    fifo_csv_dumper_772 = new("./depth772.csv");
    cstatus_csv_dumper_772 = new("./chan_status772.csv");
    fifo_monitor_772 = new(fifo_csv_dumper_772,fifo_intf_772,cstatus_csv_dumper_772);
    fifo_csv_dumper_773 = new("./depth773.csv");
    cstatus_csv_dumper_773 = new("./chan_status773.csv");
    fifo_monitor_773 = new(fifo_csv_dumper_773,fifo_intf_773,cstatus_csv_dumper_773);
    fifo_csv_dumper_774 = new("./depth774.csv");
    cstatus_csv_dumper_774 = new("./chan_status774.csv");
    fifo_monitor_774 = new(fifo_csv_dumper_774,fifo_intf_774,cstatus_csv_dumper_774);
    fifo_csv_dumper_775 = new("./depth775.csv");
    cstatus_csv_dumper_775 = new("./chan_status775.csv");
    fifo_monitor_775 = new(fifo_csv_dumper_775,fifo_intf_775,cstatus_csv_dumper_775);
    fifo_csv_dumper_776 = new("./depth776.csv");
    cstatus_csv_dumper_776 = new("./chan_status776.csv");
    fifo_monitor_776 = new(fifo_csv_dumper_776,fifo_intf_776,cstatus_csv_dumper_776);
    fifo_csv_dumper_777 = new("./depth777.csv");
    cstatus_csv_dumper_777 = new("./chan_status777.csv");
    fifo_monitor_777 = new(fifo_csv_dumper_777,fifo_intf_777,cstatus_csv_dumper_777);
    fifo_csv_dumper_778 = new("./depth778.csv");
    cstatus_csv_dumper_778 = new("./chan_status778.csv");
    fifo_monitor_778 = new(fifo_csv_dumper_778,fifo_intf_778,cstatus_csv_dumper_778);
    fifo_csv_dumper_779 = new("./depth779.csv");
    cstatus_csv_dumper_779 = new("./chan_status779.csv");
    fifo_monitor_779 = new(fifo_csv_dumper_779,fifo_intf_779,cstatus_csv_dumper_779);
    fifo_csv_dumper_780 = new("./depth780.csv");
    cstatus_csv_dumper_780 = new("./chan_status780.csv");
    fifo_monitor_780 = new(fifo_csv_dumper_780,fifo_intf_780,cstatus_csv_dumper_780);
    fifo_csv_dumper_781 = new("./depth781.csv");
    cstatus_csv_dumper_781 = new("./chan_status781.csv");
    fifo_monitor_781 = new(fifo_csv_dumper_781,fifo_intf_781,cstatus_csv_dumper_781);
    fifo_csv_dumper_782 = new("./depth782.csv");
    cstatus_csv_dumper_782 = new("./chan_status782.csv");
    fifo_monitor_782 = new(fifo_csv_dumper_782,fifo_intf_782,cstatus_csv_dumper_782);
    fifo_csv_dumper_783 = new("./depth783.csv");
    cstatus_csv_dumper_783 = new("./chan_status783.csv");
    fifo_monitor_783 = new(fifo_csv_dumper_783,fifo_intf_783,cstatus_csv_dumper_783);
    fifo_csv_dumper_784 = new("./depth784.csv");
    cstatus_csv_dumper_784 = new("./chan_status784.csv");
    fifo_monitor_784 = new(fifo_csv_dumper_784,fifo_intf_784,cstatus_csv_dumper_784);
    fifo_csv_dumper_785 = new("./depth785.csv");
    cstatus_csv_dumper_785 = new("./chan_status785.csv");
    fifo_monitor_785 = new(fifo_csv_dumper_785,fifo_intf_785,cstatus_csv_dumper_785);
    fifo_csv_dumper_786 = new("./depth786.csv");
    cstatus_csv_dumper_786 = new("./chan_status786.csv");
    fifo_monitor_786 = new(fifo_csv_dumper_786,fifo_intf_786,cstatus_csv_dumper_786);
    fifo_csv_dumper_787 = new("./depth787.csv");
    cstatus_csv_dumper_787 = new("./chan_status787.csv");
    fifo_monitor_787 = new(fifo_csv_dumper_787,fifo_intf_787,cstatus_csv_dumper_787);
    fifo_csv_dumper_788 = new("./depth788.csv");
    cstatus_csv_dumper_788 = new("./chan_status788.csv");
    fifo_monitor_788 = new(fifo_csv_dumper_788,fifo_intf_788,cstatus_csv_dumper_788);
    fifo_csv_dumper_789 = new("./depth789.csv");
    cstatus_csv_dumper_789 = new("./chan_status789.csv");
    fifo_monitor_789 = new(fifo_csv_dumper_789,fifo_intf_789,cstatus_csv_dumper_789);
    fifo_csv_dumper_790 = new("./depth790.csv");
    cstatus_csv_dumper_790 = new("./chan_status790.csv");
    fifo_monitor_790 = new(fifo_csv_dumper_790,fifo_intf_790,cstatus_csv_dumper_790);
    fifo_csv_dumper_791 = new("./depth791.csv");
    cstatus_csv_dumper_791 = new("./chan_status791.csv");
    fifo_monitor_791 = new(fifo_csv_dumper_791,fifo_intf_791,cstatus_csv_dumper_791);
    fifo_csv_dumper_792 = new("./depth792.csv");
    cstatus_csv_dumper_792 = new("./chan_status792.csv");
    fifo_monitor_792 = new(fifo_csv_dumper_792,fifo_intf_792,cstatus_csv_dumper_792);
    fifo_csv_dumper_793 = new("./depth793.csv");
    cstatus_csv_dumper_793 = new("./chan_status793.csv");
    fifo_monitor_793 = new(fifo_csv_dumper_793,fifo_intf_793,cstatus_csv_dumper_793);
    fifo_csv_dumper_794 = new("./depth794.csv");
    cstatus_csv_dumper_794 = new("./chan_status794.csv");
    fifo_monitor_794 = new(fifo_csv_dumper_794,fifo_intf_794,cstatus_csv_dumper_794);
    fifo_csv_dumper_795 = new("./depth795.csv");
    cstatus_csv_dumper_795 = new("./chan_status795.csv");
    fifo_monitor_795 = new(fifo_csv_dumper_795,fifo_intf_795,cstatus_csv_dumper_795);
    fifo_csv_dumper_796 = new("./depth796.csv");
    cstatus_csv_dumper_796 = new("./chan_status796.csv");
    fifo_monitor_796 = new(fifo_csv_dumper_796,fifo_intf_796,cstatus_csv_dumper_796);
    fifo_csv_dumper_797 = new("./depth797.csv");
    cstatus_csv_dumper_797 = new("./chan_status797.csv");
    fifo_monitor_797 = new(fifo_csv_dumper_797,fifo_intf_797,cstatus_csv_dumper_797);
    fifo_csv_dumper_798 = new("./depth798.csv");
    cstatus_csv_dumper_798 = new("./chan_status798.csv");
    fifo_monitor_798 = new(fifo_csv_dumper_798,fifo_intf_798,cstatus_csv_dumper_798);
    fifo_csv_dumper_799 = new("./depth799.csv");
    cstatus_csv_dumper_799 = new("./chan_status799.csv");
    fifo_monitor_799 = new(fifo_csv_dumper_799,fifo_intf_799,cstatus_csv_dumper_799);
    fifo_csv_dumper_800 = new("./depth800.csv");
    cstatus_csv_dumper_800 = new("./chan_status800.csv");
    fifo_monitor_800 = new(fifo_csv_dumper_800,fifo_intf_800,cstatus_csv_dumper_800);
    fifo_csv_dumper_801 = new("./depth801.csv");
    cstatus_csv_dumper_801 = new("./chan_status801.csv");
    fifo_monitor_801 = new(fifo_csv_dumper_801,fifo_intf_801,cstatus_csv_dumper_801);
    fifo_csv_dumper_802 = new("./depth802.csv");
    cstatus_csv_dumper_802 = new("./chan_status802.csv");
    fifo_monitor_802 = new(fifo_csv_dumper_802,fifo_intf_802,cstatus_csv_dumper_802);
    fifo_csv_dumper_803 = new("./depth803.csv");
    cstatus_csv_dumper_803 = new("./chan_status803.csv");
    fifo_monitor_803 = new(fifo_csv_dumper_803,fifo_intf_803,cstatus_csv_dumper_803);
    fifo_csv_dumper_804 = new("./depth804.csv");
    cstatus_csv_dumper_804 = new("./chan_status804.csv");
    fifo_monitor_804 = new(fifo_csv_dumper_804,fifo_intf_804,cstatus_csv_dumper_804);
    fifo_csv_dumper_805 = new("./depth805.csv");
    cstatus_csv_dumper_805 = new("./chan_status805.csv");
    fifo_monitor_805 = new(fifo_csv_dumper_805,fifo_intf_805,cstatus_csv_dumper_805);
    fifo_csv_dumper_806 = new("./depth806.csv");
    cstatus_csv_dumper_806 = new("./chan_status806.csv");
    fifo_monitor_806 = new(fifo_csv_dumper_806,fifo_intf_806,cstatus_csv_dumper_806);
    fifo_csv_dumper_807 = new("./depth807.csv");
    cstatus_csv_dumper_807 = new("./chan_status807.csv");
    fifo_monitor_807 = new(fifo_csv_dumper_807,fifo_intf_807,cstatus_csv_dumper_807);
    fifo_csv_dumper_808 = new("./depth808.csv");
    cstatus_csv_dumper_808 = new("./chan_status808.csv");
    fifo_monitor_808 = new(fifo_csv_dumper_808,fifo_intf_808,cstatus_csv_dumper_808);
    fifo_csv_dumper_809 = new("./depth809.csv");
    cstatus_csv_dumper_809 = new("./chan_status809.csv");
    fifo_monitor_809 = new(fifo_csv_dumper_809,fifo_intf_809,cstatus_csv_dumper_809);
    fifo_csv_dumper_810 = new("./depth810.csv");
    cstatus_csv_dumper_810 = new("./chan_status810.csv");
    fifo_monitor_810 = new(fifo_csv_dumper_810,fifo_intf_810,cstatus_csv_dumper_810);
    fifo_csv_dumper_811 = new("./depth811.csv");
    cstatus_csv_dumper_811 = new("./chan_status811.csv");
    fifo_monitor_811 = new(fifo_csv_dumper_811,fifo_intf_811,cstatus_csv_dumper_811);
    fifo_csv_dumper_812 = new("./depth812.csv");
    cstatus_csv_dumper_812 = new("./chan_status812.csv");
    fifo_monitor_812 = new(fifo_csv_dumper_812,fifo_intf_812,cstatus_csv_dumper_812);
    fifo_csv_dumper_813 = new("./depth813.csv");
    cstatus_csv_dumper_813 = new("./chan_status813.csv");
    fifo_monitor_813 = new(fifo_csv_dumper_813,fifo_intf_813,cstatus_csv_dumper_813);
    fifo_csv_dumper_814 = new("./depth814.csv");
    cstatus_csv_dumper_814 = new("./chan_status814.csv");
    fifo_monitor_814 = new(fifo_csv_dumper_814,fifo_intf_814,cstatus_csv_dumper_814);
    fifo_csv_dumper_815 = new("./depth815.csv");
    cstatus_csv_dumper_815 = new("./chan_status815.csv");
    fifo_monitor_815 = new(fifo_csv_dumper_815,fifo_intf_815,cstatus_csv_dumper_815);
    fifo_csv_dumper_816 = new("./depth816.csv");
    cstatus_csv_dumper_816 = new("./chan_status816.csv");
    fifo_monitor_816 = new(fifo_csv_dumper_816,fifo_intf_816,cstatus_csv_dumper_816);
    fifo_csv_dumper_817 = new("./depth817.csv");
    cstatus_csv_dumper_817 = new("./chan_status817.csv");
    fifo_monitor_817 = new(fifo_csv_dumper_817,fifo_intf_817,cstatus_csv_dumper_817);
    fifo_csv_dumper_818 = new("./depth818.csv");
    cstatus_csv_dumper_818 = new("./chan_status818.csv");
    fifo_monitor_818 = new(fifo_csv_dumper_818,fifo_intf_818,cstatus_csv_dumper_818);
    fifo_csv_dumper_819 = new("./depth819.csv");
    cstatus_csv_dumper_819 = new("./chan_status819.csv");
    fifo_monitor_819 = new(fifo_csv_dumper_819,fifo_intf_819,cstatus_csv_dumper_819);
    fifo_csv_dumper_820 = new("./depth820.csv");
    cstatus_csv_dumper_820 = new("./chan_status820.csv");
    fifo_monitor_820 = new(fifo_csv_dumper_820,fifo_intf_820,cstatus_csv_dumper_820);
    fifo_csv_dumper_821 = new("./depth821.csv");
    cstatus_csv_dumper_821 = new("./chan_status821.csv");
    fifo_monitor_821 = new(fifo_csv_dumper_821,fifo_intf_821,cstatus_csv_dumper_821);
    fifo_csv_dumper_822 = new("./depth822.csv");
    cstatus_csv_dumper_822 = new("./chan_status822.csv");
    fifo_monitor_822 = new(fifo_csv_dumper_822,fifo_intf_822,cstatus_csv_dumper_822);
    fifo_csv_dumper_823 = new("./depth823.csv");
    cstatus_csv_dumper_823 = new("./chan_status823.csv");
    fifo_monitor_823 = new(fifo_csv_dumper_823,fifo_intf_823,cstatus_csv_dumper_823);
    fifo_csv_dumper_824 = new("./depth824.csv");
    cstatus_csv_dumper_824 = new("./chan_status824.csv");
    fifo_monitor_824 = new(fifo_csv_dumper_824,fifo_intf_824,cstatus_csv_dumper_824);
    fifo_csv_dumper_825 = new("./depth825.csv");
    cstatus_csv_dumper_825 = new("./chan_status825.csv");
    fifo_monitor_825 = new(fifo_csv_dumper_825,fifo_intf_825,cstatus_csv_dumper_825);
    fifo_csv_dumper_826 = new("./depth826.csv");
    cstatus_csv_dumper_826 = new("./chan_status826.csv");
    fifo_monitor_826 = new(fifo_csv_dumper_826,fifo_intf_826,cstatus_csv_dumper_826);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);
    pstall_csv_dumper_6 = new("./stalling6.csv");
    pstatus_csv_dumper_6 = new("./status6.csv");
    process_monitor_6 = new(pstall_csv_dumper_6,process_intf_6,pstatus_csv_dumper_6);
    pstall_csv_dumper_7 = new("./stalling7.csv");
    pstatus_csv_dumper_7 = new("./status7.csv");
    process_monitor_7 = new(pstall_csv_dumper_7,process_intf_7,pstatus_csv_dumper_7);
    pstall_csv_dumper_8 = new("./stalling8.csv");
    pstatus_csv_dumper_8 = new("./status8.csv");
    process_monitor_8 = new(pstall_csv_dumper_8,process_intf_8,pstatus_csv_dumper_8);
    pstall_csv_dumper_9 = new("./stalling9.csv");
    pstatus_csv_dumper_9 = new("./status9.csv");
    process_monitor_9 = new(pstall_csv_dumper_9,process_intf_9,pstatus_csv_dumper_9);
    pstall_csv_dumper_10 = new("./stalling10.csv");
    pstatus_csv_dumper_10 = new("./status10.csv");
    process_monitor_10 = new(pstall_csv_dumper_10,process_intf_10,pstatus_csv_dumper_10);
    pstall_csv_dumper_11 = new("./stalling11.csv");
    pstatus_csv_dumper_11 = new("./status11.csv");
    process_monitor_11 = new(pstall_csv_dumper_11,process_intf_11,pstatus_csv_dumper_11);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);





    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(fifo_monitor_35);
    sample_manager_inst.add_one_monitor(fifo_monitor_36);
    sample_manager_inst.add_one_monitor(fifo_monitor_37);
    sample_manager_inst.add_one_monitor(fifo_monitor_38);
    sample_manager_inst.add_one_monitor(fifo_monitor_39);
    sample_manager_inst.add_one_monitor(fifo_monitor_40);
    sample_manager_inst.add_one_monitor(fifo_monitor_41);
    sample_manager_inst.add_one_monitor(fifo_monitor_42);
    sample_manager_inst.add_one_monitor(fifo_monitor_43);
    sample_manager_inst.add_one_monitor(fifo_monitor_44);
    sample_manager_inst.add_one_monitor(fifo_monitor_45);
    sample_manager_inst.add_one_monitor(fifo_monitor_46);
    sample_manager_inst.add_one_monitor(fifo_monitor_47);
    sample_manager_inst.add_one_monitor(fifo_monitor_48);
    sample_manager_inst.add_one_monitor(fifo_monitor_49);
    sample_manager_inst.add_one_monitor(fifo_monitor_50);
    sample_manager_inst.add_one_monitor(fifo_monitor_51);
    sample_manager_inst.add_one_monitor(fifo_monitor_52);
    sample_manager_inst.add_one_monitor(fifo_monitor_53);
    sample_manager_inst.add_one_monitor(fifo_monitor_54);
    sample_manager_inst.add_one_monitor(fifo_monitor_55);
    sample_manager_inst.add_one_monitor(fifo_monitor_56);
    sample_manager_inst.add_one_monitor(fifo_monitor_57);
    sample_manager_inst.add_one_monitor(fifo_monitor_58);
    sample_manager_inst.add_one_monitor(fifo_monitor_59);
    sample_manager_inst.add_one_monitor(fifo_monitor_60);
    sample_manager_inst.add_one_monitor(fifo_monitor_61);
    sample_manager_inst.add_one_monitor(fifo_monitor_62);
    sample_manager_inst.add_one_monitor(fifo_monitor_63);
    sample_manager_inst.add_one_monitor(fifo_monitor_64);
    sample_manager_inst.add_one_monitor(fifo_monitor_65);
    sample_manager_inst.add_one_monitor(fifo_monitor_66);
    sample_manager_inst.add_one_monitor(fifo_monitor_67);
    sample_manager_inst.add_one_monitor(fifo_monitor_68);
    sample_manager_inst.add_one_monitor(fifo_monitor_69);
    sample_manager_inst.add_one_monitor(fifo_monitor_70);
    sample_manager_inst.add_one_monitor(fifo_monitor_71);
    sample_manager_inst.add_one_monitor(fifo_monitor_72);
    sample_manager_inst.add_one_monitor(fifo_monitor_73);
    sample_manager_inst.add_one_monitor(fifo_monitor_74);
    sample_manager_inst.add_one_monitor(fifo_monitor_75);
    sample_manager_inst.add_one_monitor(fifo_monitor_76);
    sample_manager_inst.add_one_monitor(fifo_monitor_77);
    sample_manager_inst.add_one_monitor(fifo_monitor_78);
    sample_manager_inst.add_one_monitor(fifo_monitor_79);
    sample_manager_inst.add_one_monitor(fifo_monitor_80);
    sample_manager_inst.add_one_monitor(fifo_monitor_81);
    sample_manager_inst.add_one_monitor(fifo_monitor_82);
    sample_manager_inst.add_one_monitor(fifo_monitor_83);
    sample_manager_inst.add_one_monitor(fifo_monitor_84);
    sample_manager_inst.add_one_monitor(fifo_monitor_85);
    sample_manager_inst.add_one_monitor(fifo_monitor_86);
    sample_manager_inst.add_one_monitor(fifo_monitor_87);
    sample_manager_inst.add_one_monitor(fifo_monitor_88);
    sample_manager_inst.add_one_monitor(fifo_monitor_89);
    sample_manager_inst.add_one_monitor(fifo_monitor_90);
    sample_manager_inst.add_one_monitor(fifo_monitor_91);
    sample_manager_inst.add_one_monitor(fifo_monitor_92);
    sample_manager_inst.add_one_monitor(fifo_monitor_93);
    sample_manager_inst.add_one_monitor(fifo_monitor_94);
    sample_manager_inst.add_one_monitor(fifo_monitor_95);
    sample_manager_inst.add_one_monitor(fifo_monitor_96);
    sample_manager_inst.add_one_monitor(fifo_monitor_97);
    sample_manager_inst.add_one_monitor(fifo_monitor_98);
    sample_manager_inst.add_one_monitor(fifo_monitor_99);
    sample_manager_inst.add_one_monitor(fifo_monitor_100);
    sample_manager_inst.add_one_monitor(fifo_monitor_101);
    sample_manager_inst.add_one_monitor(fifo_monitor_102);
    sample_manager_inst.add_one_monitor(fifo_monitor_103);
    sample_manager_inst.add_one_monitor(fifo_monitor_104);
    sample_manager_inst.add_one_monitor(fifo_monitor_105);
    sample_manager_inst.add_one_monitor(fifo_monitor_106);
    sample_manager_inst.add_one_monitor(fifo_monitor_107);
    sample_manager_inst.add_one_monitor(fifo_monitor_108);
    sample_manager_inst.add_one_monitor(fifo_monitor_109);
    sample_manager_inst.add_one_monitor(fifo_monitor_110);
    sample_manager_inst.add_one_monitor(fifo_monitor_111);
    sample_manager_inst.add_one_monitor(fifo_monitor_112);
    sample_manager_inst.add_one_monitor(fifo_monitor_113);
    sample_manager_inst.add_one_monitor(fifo_monitor_114);
    sample_manager_inst.add_one_monitor(fifo_monitor_115);
    sample_manager_inst.add_one_monitor(fifo_monitor_116);
    sample_manager_inst.add_one_monitor(fifo_monitor_117);
    sample_manager_inst.add_one_monitor(fifo_monitor_118);
    sample_manager_inst.add_one_monitor(fifo_monitor_119);
    sample_manager_inst.add_one_monitor(fifo_monitor_120);
    sample_manager_inst.add_one_monitor(fifo_monitor_121);
    sample_manager_inst.add_one_monitor(fifo_monitor_122);
    sample_manager_inst.add_one_monitor(fifo_monitor_123);
    sample_manager_inst.add_one_monitor(fifo_monitor_124);
    sample_manager_inst.add_one_monitor(fifo_monitor_125);
    sample_manager_inst.add_one_monitor(fifo_monitor_126);
    sample_manager_inst.add_one_monitor(fifo_monitor_127);
    sample_manager_inst.add_one_monitor(fifo_monitor_128);
    sample_manager_inst.add_one_monitor(fifo_monitor_129);
    sample_manager_inst.add_one_monitor(fifo_monitor_130);
    sample_manager_inst.add_one_monitor(fifo_monitor_131);
    sample_manager_inst.add_one_monitor(fifo_monitor_132);
    sample_manager_inst.add_one_monitor(fifo_monitor_133);
    sample_manager_inst.add_one_monitor(fifo_monitor_134);
    sample_manager_inst.add_one_monitor(fifo_monitor_135);
    sample_manager_inst.add_one_monitor(fifo_monitor_136);
    sample_manager_inst.add_one_monitor(fifo_monitor_137);
    sample_manager_inst.add_one_monitor(fifo_monitor_138);
    sample_manager_inst.add_one_monitor(fifo_monitor_139);
    sample_manager_inst.add_one_monitor(fifo_monitor_140);
    sample_manager_inst.add_one_monitor(fifo_monitor_141);
    sample_manager_inst.add_one_monitor(fifo_monitor_142);
    sample_manager_inst.add_one_monitor(fifo_monitor_143);
    sample_manager_inst.add_one_monitor(fifo_monitor_144);
    sample_manager_inst.add_one_monitor(fifo_monitor_145);
    sample_manager_inst.add_one_monitor(fifo_monitor_146);
    sample_manager_inst.add_one_monitor(fifo_monitor_147);
    sample_manager_inst.add_one_monitor(fifo_monitor_148);
    sample_manager_inst.add_one_monitor(fifo_monitor_149);
    sample_manager_inst.add_one_monitor(fifo_monitor_150);
    sample_manager_inst.add_one_monitor(fifo_monitor_151);
    sample_manager_inst.add_one_monitor(fifo_monitor_152);
    sample_manager_inst.add_one_monitor(fifo_monitor_153);
    sample_manager_inst.add_one_monitor(fifo_monitor_154);
    sample_manager_inst.add_one_monitor(fifo_monitor_155);
    sample_manager_inst.add_one_monitor(fifo_monitor_156);
    sample_manager_inst.add_one_monitor(fifo_monitor_157);
    sample_manager_inst.add_one_monitor(fifo_monitor_158);
    sample_manager_inst.add_one_monitor(fifo_monitor_159);
    sample_manager_inst.add_one_monitor(fifo_monitor_160);
    sample_manager_inst.add_one_monitor(fifo_monitor_161);
    sample_manager_inst.add_one_monitor(fifo_monitor_162);
    sample_manager_inst.add_one_monitor(fifo_monitor_163);
    sample_manager_inst.add_one_monitor(fifo_monitor_164);
    sample_manager_inst.add_one_monitor(fifo_monitor_165);
    sample_manager_inst.add_one_monitor(fifo_monitor_166);
    sample_manager_inst.add_one_monitor(fifo_monitor_167);
    sample_manager_inst.add_one_monitor(fifo_monitor_168);
    sample_manager_inst.add_one_monitor(fifo_monitor_169);
    sample_manager_inst.add_one_monitor(fifo_monitor_170);
    sample_manager_inst.add_one_monitor(fifo_monitor_171);
    sample_manager_inst.add_one_monitor(fifo_monitor_172);
    sample_manager_inst.add_one_monitor(fifo_monitor_173);
    sample_manager_inst.add_one_monitor(fifo_monitor_174);
    sample_manager_inst.add_one_monitor(fifo_monitor_175);
    sample_manager_inst.add_one_monitor(fifo_monitor_176);
    sample_manager_inst.add_one_monitor(fifo_monitor_177);
    sample_manager_inst.add_one_monitor(fifo_monitor_178);
    sample_manager_inst.add_one_monitor(fifo_monitor_179);
    sample_manager_inst.add_one_monitor(fifo_monitor_180);
    sample_manager_inst.add_one_monitor(fifo_monitor_181);
    sample_manager_inst.add_one_monitor(fifo_monitor_182);
    sample_manager_inst.add_one_monitor(fifo_monitor_183);
    sample_manager_inst.add_one_monitor(fifo_monitor_184);
    sample_manager_inst.add_one_monitor(fifo_monitor_185);
    sample_manager_inst.add_one_monitor(fifo_monitor_186);
    sample_manager_inst.add_one_monitor(fifo_monitor_187);
    sample_manager_inst.add_one_monitor(fifo_monitor_188);
    sample_manager_inst.add_one_monitor(fifo_monitor_189);
    sample_manager_inst.add_one_monitor(fifo_monitor_190);
    sample_manager_inst.add_one_monitor(fifo_monitor_191);
    sample_manager_inst.add_one_monitor(fifo_monitor_192);
    sample_manager_inst.add_one_monitor(fifo_monitor_193);
    sample_manager_inst.add_one_monitor(fifo_monitor_194);
    sample_manager_inst.add_one_monitor(fifo_monitor_195);
    sample_manager_inst.add_one_monitor(fifo_monitor_196);
    sample_manager_inst.add_one_monitor(fifo_monitor_197);
    sample_manager_inst.add_one_monitor(fifo_monitor_198);
    sample_manager_inst.add_one_monitor(fifo_monitor_199);
    sample_manager_inst.add_one_monitor(fifo_monitor_200);
    sample_manager_inst.add_one_monitor(fifo_monitor_201);
    sample_manager_inst.add_one_monitor(fifo_monitor_202);
    sample_manager_inst.add_one_monitor(fifo_monitor_203);
    sample_manager_inst.add_one_monitor(fifo_monitor_204);
    sample_manager_inst.add_one_monitor(fifo_monitor_205);
    sample_manager_inst.add_one_monitor(fifo_monitor_206);
    sample_manager_inst.add_one_monitor(fifo_monitor_207);
    sample_manager_inst.add_one_monitor(fifo_monitor_208);
    sample_manager_inst.add_one_monitor(fifo_monitor_209);
    sample_manager_inst.add_one_monitor(fifo_monitor_210);
    sample_manager_inst.add_one_monitor(fifo_monitor_211);
    sample_manager_inst.add_one_monitor(fifo_monitor_212);
    sample_manager_inst.add_one_monitor(fifo_monitor_213);
    sample_manager_inst.add_one_monitor(fifo_monitor_214);
    sample_manager_inst.add_one_monitor(fifo_monitor_215);
    sample_manager_inst.add_one_monitor(fifo_monitor_216);
    sample_manager_inst.add_one_monitor(fifo_monitor_217);
    sample_manager_inst.add_one_monitor(fifo_monitor_218);
    sample_manager_inst.add_one_monitor(fifo_monitor_219);
    sample_manager_inst.add_one_monitor(fifo_monitor_220);
    sample_manager_inst.add_one_monitor(fifo_monitor_221);
    sample_manager_inst.add_one_monitor(fifo_monitor_222);
    sample_manager_inst.add_one_monitor(fifo_monitor_223);
    sample_manager_inst.add_one_monitor(fifo_monitor_224);
    sample_manager_inst.add_one_monitor(fifo_monitor_225);
    sample_manager_inst.add_one_monitor(fifo_monitor_226);
    sample_manager_inst.add_one_monitor(fifo_monitor_227);
    sample_manager_inst.add_one_monitor(fifo_monitor_228);
    sample_manager_inst.add_one_monitor(fifo_monitor_229);
    sample_manager_inst.add_one_monitor(fifo_monitor_230);
    sample_manager_inst.add_one_monitor(fifo_monitor_231);
    sample_manager_inst.add_one_monitor(fifo_monitor_232);
    sample_manager_inst.add_one_monitor(fifo_monitor_233);
    sample_manager_inst.add_one_monitor(fifo_monitor_234);
    sample_manager_inst.add_one_monitor(fifo_monitor_235);
    sample_manager_inst.add_one_monitor(fifo_monitor_236);
    sample_manager_inst.add_one_monitor(fifo_monitor_237);
    sample_manager_inst.add_one_monitor(fifo_monitor_238);
    sample_manager_inst.add_one_monitor(fifo_monitor_239);
    sample_manager_inst.add_one_monitor(fifo_monitor_240);
    sample_manager_inst.add_one_monitor(fifo_monitor_241);
    sample_manager_inst.add_one_monitor(fifo_monitor_242);
    sample_manager_inst.add_one_monitor(fifo_monitor_243);
    sample_manager_inst.add_one_monitor(fifo_monitor_244);
    sample_manager_inst.add_one_monitor(fifo_monitor_245);
    sample_manager_inst.add_one_monitor(fifo_monitor_246);
    sample_manager_inst.add_one_monitor(fifo_monitor_247);
    sample_manager_inst.add_one_monitor(fifo_monitor_248);
    sample_manager_inst.add_one_monitor(fifo_monitor_249);
    sample_manager_inst.add_one_monitor(fifo_monitor_250);
    sample_manager_inst.add_one_monitor(fifo_monitor_251);
    sample_manager_inst.add_one_monitor(fifo_monitor_252);
    sample_manager_inst.add_one_monitor(fifo_monitor_253);
    sample_manager_inst.add_one_monitor(fifo_monitor_254);
    sample_manager_inst.add_one_monitor(fifo_monitor_255);
    sample_manager_inst.add_one_monitor(fifo_monitor_256);
    sample_manager_inst.add_one_monitor(fifo_monitor_257);
    sample_manager_inst.add_one_monitor(fifo_monitor_258);
    sample_manager_inst.add_one_monitor(fifo_monitor_259);
    sample_manager_inst.add_one_monitor(fifo_monitor_260);
    sample_manager_inst.add_one_monitor(fifo_monitor_261);
    sample_manager_inst.add_one_monitor(fifo_monitor_262);
    sample_manager_inst.add_one_monitor(fifo_monitor_263);
    sample_manager_inst.add_one_monitor(fifo_monitor_264);
    sample_manager_inst.add_one_monitor(fifo_monitor_265);
    sample_manager_inst.add_one_monitor(fifo_monitor_266);
    sample_manager_inst.add_one_monitor(fifo_monitor_267);
    sample_manager_inst.add_one_monitor(fifo_monitor_268);
    sample_manager_inst.add_one_monitor(fifo_monitor_269);
    sample_manager_inst.add_one_monitor(fifo_monitor_270);
    sample_manager_inst.add_one_monitor(fifo_monitor_271);
    sample_manager_inst.add_one_monitor(fifo_monitor_272);
    sample_manager_inst.add_one_monitor(fifo_monitor_273);
    sample_manager_inst.add_one_monitor(fifo_monitor_274);
    sample_manager_inst.add_one_monitor(fifo_monitor_275);
    sample_manager_inst.add_one_monitor(fifo_monitor_276);
    sample_manager_inst.add_one_monitor(fifo_monitor_277);
    sample_manager_inst.add_one_monitor(fifo_monitor_278);
    sample_manager_inst.add_one_monitor(fifo_monitor_279);
    sample_manager_inst.add_one_monitor(fifo_monitor_280);
    sample_manager_inst.add_one_monitor(fifo_monitor_281);
    sample_manager_inst.add_one_monitor(fifo_monitor_282);
    sample_manager_inst.add_one_monitor(fifo_monitor_283);
    sample_manager_inst.add_one_monitor(fifo_monitor_284);
    sample_manager_inst.add_one_monitor(fifo_monitor_285);
    sample_manager_inst.add_one_monitor(fifo_monitor_286);
    sample_manager_inst.add_one_monitor(fifo_monitor_287);
    sample_manager_inst.add_one_monitor(fifo_monitor_288);
    sample_manager_inst.add_one_monitor(fifo_monitor_289);
    sample_manager_inst.add_one_monitor(fifo_monitor_290);
    sample_manager_inst.add_one_monitor(fifo_monitor_291);
    sample_manager_inst.add_one_monitor(fifo_monitor_292);
    sample_manager_inst.add_one_monitor(fifo_monitor_293);
    sample_manager_inst.add_one_monitor(fifo_monitor_294);
    sample_manager_inst.add_one_monitor(fifo_monitor_295);
    sample_manager_inst.add_one_monitor(fifo_monitor_296);
    sample_manager_inst.add_one_monitor(fifo_monitor_297);
    sample_manager_inst.add_one_monitor(fifo_monitor_298);
    sample_manager_inst.add_one_monitor(fifo_monitor_299);
    sample_manager_inst.add_one_monitor(fifo_monitor_300);
    sample_manager_inst.add_one_monitor(fifo_monitor_301);
    sample_manager_inst.add_one_monitor(fifo_monitor_302);
    sample_manager_inst.add_one_monitor(fifo_monitor_303);
    sample_manager_inst.add_one_monitor(fifo_monitor_304);
    sample_manager_inst.add_one_monitor(fifo_monitor_305);
    sample_manager_inst.add_one_monitor(fifo_monitor_306);
    sample_manager_inst.add_one_monitor(fifo_monitor_307);
    sample_manager_inst.add_one_monitor(fifo_monitor_308);
    sample_manager_inst.add_one_monitor(fifo_monitor_309);
    sample_manager_inst.add_one_monitor(fifo_monitor_310);
    sample_manager_inst.add_one_monitor(fifo_monitor_311);
    sample_manager_inst.add_one_monitor(fifo_monitor_312);
    sample_manager_inst.add_one_monitor(fifo_monitor_313);
    sample_manager_inst.add_one_monitor(fifo_monitor_314);
    sample_manager_inst.add_one_monitor(fifo_monitor_315);
    sample_manager_inst.add_one_monitor(fifo_monitor_316);
    sample_manager_inst.add_one_monitor(fifo_monitor_317);
    sample_manager_inst.add_one_monitor(fifo_monitor_318);
    sample_manager_inst.add_one_monitor(fifo_monitor_319);
    sample_manager_inst.add_one_monitor(fifo_monitor_320);
    sample_manager_inst.add_one_monitor(fifo_monitor_321);
    sample_manager_inst.add_one_monitor(fifo_monitor_322);
    sample_manager_inst.add_one_monitor(fifo_monitor_323);
    sample_manager_inst.add_one_monitor(fifo_monitor_324);
    sample_manager_inst.add_one_monitor(fifo_monitor_325);
    sample_manager_inst.add_one_monitor(fifo_monitor_326);
    sample_manager_inst.add_one_monitor(fifo_monitor_327);
    sample_manager_inst.add_one_monitor(fifo_monitor_328);
    sample_manager_inst.add_one_monitor(fifo_monitor_329);
    sample_manager_inst.add_one_monitor(fifo_monitor_330);
    sample_manager_inst.add_one_monitor(fifo_monitor_331);
    sample_manager_inst.add_one_monitor(fifo_monitor_332);
    sample_manager_inst.add_one_monitor(fifo_monitor_333);
    sample_manager_inst.add_one_monitor(fifo_monitor_334);
    sample_manager_inst.add_one_monitor(fifo_monitor_335);
    sample_manager_inst.add_one_monitor(fifo_monitor_336);
    sample_manager_inst.add_one_monitor(fifo_monitor_337);
    sample_manager_inst.add_one_monitor(fifo_monitor_338);
    sample_manager_inst.add_one_monitor(fifo_monitor_339);
    sample_manager_inst.add_one_monitor(fifo_monitor_340);
    sample_manager_inst.add_one_monitor(fifo_monitor_341);
    sample_manager_inst.add_one_monitor(fifo_monitor_342);
    sample_manager_inst.add_one_monitor(fifo_monitor_343);
    sample_manager_inst.add_one_monitor(fifo_monitor_344);
    sample_manager_inst.add_one_monitor(fifo_monitor_345);
    sample_manager_inst.add_one_monitor(fifo_monitor_346);
    sample_manager_inst.add_one_monitor(fifo_monitor_347);
    sample_manager_inst.add_one_monitor(fifo_monitor_348);
    sample_manager_inst.add_one_monitor(fifo_monitor_349);
    sample_manager_inst.add_one_monitor(fifo_monitor_350);
    sample_manager_inst.add_one_monitor(fifo_monitor_351);
    sample_manager_inst.add_one_monitor(fifo_monitor_352);
    sample_manager_inst.add_one_monitor(fifo_monitor_353);
    sample_manager_inst.add_one_monitor(fifo_monitor_354);
    sample_manager_inst.add_one_monitor(fifo_monitor_355);
    sample_manager_inst.add_one_monitor(fifo_monitor_356);
    sample_manager_inst.add_one_monitor(fifo_monitor_357);
    sample_manager_inst.add_one_monitor(fifo_monitor_358);
    sample_manager_inst.add_one_monitor(fifo_monitor_359);
    sample_manager_inst.add_one_monitor(fifo_monitor_360);
    sample_manager_inst.add_one_monitor(fifo_monitor_361);
    sample_manager_inst.add_one_monitor(fifo_monitor_362);
    sample_manager_inst.add_one_monitor(fifo_monitor_363);
    sample_manager_inst.add_one_monitor(fifo_monitor_364);
    sample_manager_inst.add_one_monitor(fifo_monitor_365);
    sample_manager_inst.add_one_monitor(fifo_monitor_366);
    sample_manager_inst.add_one_monitor(fifo_monitor_367);
    sample_manager_inst.add_one_monitor(fifo_monitor_368);
    sample_manager_inst.add_one_monitor(fifo_monitor_369);
    sample_manager_inst.add_one_monitor(fifo_monitor_370);
    sample_manager_inst.add_one_monitor(fifo_monitor_371);
    sample_manager_inst.add_one_monitor(fifo_monitor_372);
    sample_manager_inst.add_one_monitor(fifo_monitor_373);
    sample_manager_inst.add_one_monitor(fifo_monitor_374);
    sample_manager_inst.add_one_monitor(fifo_monitor_375);
    sample_manager_inst.add_one_monitor(fifo_monitor_376);
    sample_manager_inst.add_one_monitor(fifo_monitor_377);
    sample_manager_inst.add_one_monitor(fifo_monitor_378);
    sample_manager_inst.add_one_monitor(fifo_monitor_379);
    sample_manager_inst.add_one_monitor(fifo_monitor_380);
    sample_manager_inst.add_one_monitor(fifo_monitor_381);
    sample_manager_inst.add_one_monitor(fifo_monitor_382);
    sample_manager_inst.add_one_monitor(fifo_monitor_383);
    sample_manager_inst.add_one_monitor(fifo_monitor_384);
    sample_manager_inst.add_one_monitor(fifo_monitor_385);
    sample_manager_inst.add_one_monitor(fifo_monitor_386);
    sample_manager_inst.add_one_monitor(fifo_monitor_387);
    sample_manager_inst.add_one_monitor(fifo_monitor_388);
    sample_manager_inst.add_one_monitor(fifo_monitor_389);
    sample_manager_inst.add_one_monitor(fifo_monitor_390);
    sample_manager_inst.add_one_monitor(fifo_monitor_391);
    sample_manager_inst.add_one_monitor(fifo_monitor_392);
    sample_manager_inst.add_one_monitor(fifo_monitor_393);
    sample_manager_inst.add_one_monitor(fifo_monitor_394);
    sample_manager_inst.add_one_monitor(fifo_monitor_395);
    sample_manager_inst.add_one_monitor(fifo_monitor_396);
    sample_manager_inst.add_one_monitor(fifo_monitor_397);
    sample_manager_inst.add_one_monitor(fifo_monitor_398);
    sample_manager_inst.add_one_monitor(fifo_monitor_399);
    sample_manager_inst.add_one_monitor(fifo_monitor_400);
    sample_manager_inst.add_one_monitor(fifo_monitor_401);
    sample_manager_inst.add_one_monitor(fifo_monitor_402);
    sample_manager_inst.add_one_monitor(fifo_monitor_403);
    sample_manager_inst.add_one_monitor(fifo_monitor_404);
    sample_manager_inst.add_one_monitor(fifo_monitor_405);
    sample_manager_inst.add_one_monitor(fifo_monitor_406);
    sample_manager_inst.add_one_monitor(fifo_monitor_407);
    sample_manager_inst.add_one_monitor(fifo_monitor_408);
    sample_manager_inst.add_one_monitor(fifo_monitor_409);
    sample_manager_inst.add_one_monitor(fifo_monitor_410);
    sample_manager_inst.add_one_monitor(fifo_monitor_411);
    sample_manager_inst.add_one_monitor(fifo_monitor_412);
    sample_manager_inst.add_one_monitor(fifo_monitor_413);
    sample_manager_inst.add_one_monitor(fifo_monitor_414);
    sample_manager_inst.add_one_monitor(fifo_monitor_415);
    sample_manager_inst.add_one_monitor(fifo_monitor_416);
    sample_manager_inst.add_one_monitor(fifo_monitor_417);
    sample_manager_inst.add_one_monitor(fifo_monitor_418);
    sample_manager_inst.add_one_monitor(fifo_monitor_419);
    sample_manager_inst.add_one_monitor(fifo_monitor_420);
    sample_manager_inst.add_one_monitor(fifo_monitor_421);
    sample_manager_inst.add_one_monitor(fifo_monitor_422);
    sample_manager_inst.add_one_monitor(fifo_monitor_423);
    sample_manager_inst.add_one_monitor(fifo_monitor_424);
    sample_manager_inst.add_one_monitor(fifo_monitor_425);
    sample_manager_inst.add_one_monitor(fifo_monitor_426);
    sample_manager_inst.add_one_monitor(fifo_monitor_427);
    sample_manager_inst.add_one_monitor(fifo_monitor_428);
    sample_manager_inst.add_one_monitor(fifo_monitor_429);
    sample_manager_inst.add_one_monitor(fifo_monitor_430);
    sample_manager_inst.add_one_monitor(fifo_monitor_431);
    sample_manager_inst.add_one_monitor(fifo_monitor_432);
    sample_manager_inst.add_one_monitor(fifo_monitor_433);
    sample_manager_inst.add_one_monitor(fifo_monitor_434);
    sample_manager_inst.add_one_monitor(fifo_monitor_435);
    sample_manager_inst.add_one_monitor(fifo_monitor_436);
    sample_manager_inst.add_one_monitor(fifo_monitor_437);
    sample_manager_inst.add_one_monitor(fifo_monitor_438);
    sample_manager_inst.add_one_monitor(fifo_monitor_439);
    sample_manager_inst.add_one_monitor(fifo_monitor_440);
    sample_manager_inst.add_one_monitor(fifo_monitor_441);
    sample_manager_inst.add_one_monitor(fifo_monitor_442);
    sample_manager_inst.add_one_monitor(fifo_monitor_443);
    sample_manager_inst.add_one_monitor(fifo_monitor_444);
    sample_manager_inst.add_one_monitor(fifo_monitor_445);
    sample_manager_inst.add_one_monitor(fifo_monitor_446);
    sample_manager_inst.add_one_monitor(fifo_monitor_447);
    sample_manager_inst.add_one_monitor(fifo_monitor_448);
    sample_manager_inst.add_one_monitor(fifo_monitor_449);
    sample_manager_inst.add_one_monitor(fifo_monitor_450);
    sample_manager_inst.add_one_monitor(fifo_monitor_451);
    sample_manager_inst.add_one_monitor(fifo_monitor_452);
    sample_manager_inst.add_one_monitor(fifo_monitor_453);
    sample_manager_inst.add_one_monitor(fifo_monitor_454);
    sample_manager_inst.add_one_monitor(fifo_monitor_455);
    sample_manager_inst.add_one_monitor(fifo_monitor_456);
    sample_manager_inst.add_one_monitor(fifo_monitor_457);
    sample_manager_inst.add_one_monitor(fifo_monitor_458);
    sample_manager_inst.add_one_monitor(fifo_monitor_459);
    sample_manager_inst.add_one_monitor(fifo_monitor_460);
    sample_manager_inst.add_one_monitor(fifo_monitor_461);
    sample_manager_inst.add_one_monitor(fifo_monitor_462);
    sample_manager_inst.add_one_monitor(fifo_monitor_463);
    sample_manager_inst.add_one_monitor(fifo_monitor_464);
    sample_manager_inst.add_one_monitor(fifo_monitor_465);
    sample_manager_inst.add_one_monitor(fifo_monitor_466);
    sample_manager_inst.add_one_monitor(fifo_monitor_467);
    sample_manager_inst.add_one_monitor(fifo_monitor_468);
    sample_manager_inst.add_one_monitor(fifo_monitor_469);
    sample_manager_inst.add_one_monitor(fifo_monitor_470);
    sample_manager_inst.add_one_monitor(fifo_monitor_471);
    sample_manager_inst.add_one_monitor(fifo_monitor_472);
    sample_manager_inst.add_one_monitor(fifo_monitor_473);
    sample_manager_inst.add_one_monitor(fifo_monitor_474);
    sample_manager_inst.add_one_monitor(fifo_monitor_475);
    sample_manager_inst.add_one_monitor(fifo_monitor_476);
    sample_manager_inst.add_one_monitor(fifo_monitor_477);
    sample_manager_inst.add_one_monitor(fifo_monitor_478);
    sample_manager_inst.add_one_monitor(fifo_monitor_479);
    sample_manager_inst.add_one_monitor(fifo_monitor_480);
    sample_manager_inst.add_one_monitor(fifo_monitor_481);
    sample_manager_inst.add_one_monitor(fifo_monitor_482);
    sample_manager_inst.add_one_monitor(fifo_monitor_483);
    sample_manager_inst.add_one_monitor(fifo_monitor_484);
    sample_manager_inst.add_one_monitor(fifo_monitor_485);
    sample_manager_inst.add_one_monitor(fifo_monitor_486);
    sample_manager_inst.add_one_monitor(fifo_monitor_487);
    sample_manager_inst.add_one_monitor(fifo_monitor_488);
    sample_manager_inst.add_one_monitor(fifo_monitor_489);
    sample_manager_inst.add_one_monitor(fifo_monitor_490);
    sample_manager_inst.add_one_monitor(fifo_monitor_491);
    sample_manager_inst.add_one_monitor(fifo_monitor_492);
    sample_manager_inst.add_one_monitor(fifo_monitor_493);
    sample_manager_inst.add_one_monitor(fifo_monitor_494);
    sample_manager_inst.add_one_monitor(fifo_monitor_495);
    sample_manager_inst.add_one_monitor(fifo_monitor_496);
    sample_manager_inst.add_one_monitor(fifo_monitor_497);
    sample_manager_inst.add_one_monitor(fifo_monitor_498);
    sample_manager_inst.add_one_monitor(fifo_monitor_499);
    sample_manager_inst.add_one_monitor(fifo_monitor_500);
    sample_manager_inst.add_one_monitor(fifo_monitor_501);
    sample_manager_inst.add_one_monitor(fifo_monitor_502);
    sample_manager_inst.add_one_monitor(fifo_monitor_503);
    sample_manager_inst.add_one_monitor(fifo_monitor_504);
    sample_manager_inst.add_one_monitor(fifo_monitor_505);
    sample_manager_inst.add_one_monitor(fifo_monitor_506);
    sample_manager_inst.add_one_monitor(fifo_monitor_507);
    sample_manager_inst.add_one_monitor(fifo_monitor_508);
    sample_manager_inst.add_one_monitor(fifo_monitor_509);
    sample_manager_inst.add_one_monitor(fifo_monitor_510);
    sample_manager_inst.add_one_monitor(fifo_monitor_511);
    sample_manager_inst.add_one_monitor(fifo_monitor_512);
    sample_manager_inst.add_one_monitor(fifo_monitor_513);
    sample_manager_inst.add_one_monitor(fifo_monitor_514);
    sample_manager_inst.add_one_monitor(fifo_monitor_515);
    sample_manager_inst.add_one_monitor(fifo_monitor_516);
    sample_manager_inst.add_one_monitor(fifo_monitor_517);
    sample_manager_inst.add_one_monitor(fifo_monitor_518);
    sample_manager_inst.add_one_monitor(fifo_monitor_519);
    sample_manager_inst.add_one_monitor(fifo_monitor_520);
    sample_manager_inst.add_one_monitor(fifo_monitor_521);
    sample_manager_inst.add_one_monitor(fifo_monitor_522);
    sample_manager_inst.add_one_monitor(fifo_monitor_523);
    sample_manager_inst.add_one_monitor(fifo_monitor_524);
    sample_manager_inst.add_one_monitor(fifo_monitor_525);
    sample_manager_inst.add_one_monitor(fifo_monitor_526);
    sample_manager_inst.add_one_monitor(fifo_monitor_527);
    sample_manager_inst.add_one_monitor(fifo_monitor_528);
    sample_manager_inst.add_one_monitor(fifo_monitor_529);
    sample_manager_inst.add_one_monitor(fifo_monitor_530);
    sample_manager_inst.add_one_monitor(fifo_monitor_531);
    sample_manager_inst.add_one_monitor(fifo_monitor_532);
    sample_manager_inst.add_one_monitor(fifo_monitor_533);
    sample_manager_inst.add_one_monitor(fifo_monitor_534);
    sample_manager_inst.add_one_monitor(fifo_monitor_535);
    sample_manager_inst.add_one_monitor(fifo_monitor_536);
    sample_manager_inst.add_one_monitor(fifo_monitor_537);
    sample_manager_inst.add_one_monitor(fifo_monitor_538);
    sample_manager_inst.add_one_monitor(fifo_monitor_539);
    sample_manager_inst.add_one_monitor(fifo_monitor_540);
    sample_manager_inst.add_one_monitor(fifo_monitor_541);
    sample_manager_inst.add_one_monitor(fifo_monitor_542);
    sample_manager_inst.add_one_monitor(fifo_monitor_543);
    sample_manager_inst.add_one_monitor(fifo_monitor_544);
    sample_manager_inst.add_one_monitor(fifo_monitor_545);
    sample_manager_inst.add_one_monitor(fifo_monitor_546);
    sample_manager_inst.add_one_monitor(fifo_monitor_547);
    sample_manager_inst.add_one_monitor(fifo_monitor_548);
    sample_manager_inst.add_one_monitor(fifo_monitor_549);
    sample_manager_inst.add_one_monitor(fifo_monitor_550);
    sample_manager_inst.add_one_monitor(fifo_monitor_551);
    sample_manager_inst.add_one_monitor(fifo_monitor_552);
    sample_manager_inst.add_one_monitor(fifo_monitor_553);
    sample_manager_inst.add_one_monitor(fifo_monitor_554);
    sample_manager_inst.add_one_monitor(fifo_monitor_555);
    sample_manager_inst.add_one_monitor(fifo_monitor_556);
    sample_manager_inst.add_one_monitor(fifo_monitor_557);
    sample_manager_inst.add_one_monitor(fifo_monitor_558);
    sample_manager_inst.add_one_monitor(fifo_monitor_559);
    sample_manager_inst.add_one_monitor(fifo_monitor_560);
    sample_manager_inst.add_one_monitor(fifo_monitor_561);
    sample_manager_inst.add_one_monitor(fifo_monitor_562);
    sample_manager_inst.add_one_monitor(fifo_monitor_563);
    sample_manager_inst.add_one_monitor(fifo_monitor_564);
    sample_manager_inst.add_one_monitor(fifo_monitor_565);
    sample_manager_inst.add_one_monitor(fifo_monitor_566);
    sample_manager_inst.add_one_monitor(fifo_monitor_567);
    sample_manager_inst.add_one_monitor(fifo_monitor_568);
    sample_manager_inst.add_one_monitor(fifo_monitor_569);
    sample_manager_inst.add_one_monitor(fifo_monitor_570);
    sample_manager_inst.add_one_monitor(fifo_monitor_571);
    sample_manager_inst.add_one_monitor(fifo_monitor_572);
    sample_manager_inst.add_one_monitor(fifo_monitor_573);
    sample_manager_inst.add_one_monitor(fifo_monitor_574);
    sample_manager_inst.add_one_monitor(fifo_monitor_575);
    sample_manager_inst.add_one_monitor(fifo_monitor_576);
    sample_manager_inst.add_one_monitor(fifo_monitor_577);
    sample_manager_inst.add_one_monitor(fifo_monitor_578);
    sample_manager_inst.add_one_monitor(fifo_monitor_579);
    sample_manager_inst.add_one_monitor(fifo_monitor_580);
    sample_manager_inst.add_one_monitor(fifo_monitor_581);
    sample_manager_inst.add_one_monitor(fifo_monitor_582);
    sample_manager_inst.add_one_monitor(fifo_monitor_583);
    sample_manager_inst.add_one_monitor(fifo_monitor_584);
    sample_manager_inst.add_one_monitor(fifo_monitor_585);
    sample_manager_inst.add_one_monitor(fifo_monitor_586);
    sample_manager_inst.add_one_monitor(fifo_monitor_587);
    sample_manager_inst.add_one_monitor(fifo_monitor_588);
    sample_manager_inst.add_one_monitor(fifo_monitor_589);
    sample_manager_inst.add_one_monitor(fifo_monitor_590);
    sample_manager_inst.add_one_monitor(fifo_monitor_591);
    sample_manager_inst.add_one_monitor(fifo_monitor_592);
    sample_manager_inst.add_one_monitor(fifo_monitor_593);
    sample_manager_inst.add_one_monitor(fifo_monitor_594);
    sample_manager_inst.add_one_monitor(fifo_monitor_595);
    sample_manager_inst.add_one_monitor(fifo_monitor_596);
    sample_manager_inst.add_one_monitor(fifo_monitor_597);
    sample_manager_inst.add_one_monitor(fifo_monitor_598);
    sample_manager_inst.add_one_monitor(fifo_monitor_599);
    sample_manager_inst.add_one_monitor(fifo_monitor_600);
    sample_manager_inst.add_one_monitor(fifo_monitor_601);
    sample_manager_inst.add_one_monitor(fifo_monitor_602);
    sample_manager_inst.add_one_monitor(fifo_monitor_603);
    sample_manager_inst.add_one_monitor(fifo_monitor_604);
    sample_manager_inst.add_one_monitor(fifo_monitor_605);
    sample_manager_inst.add_one_monitor(fifo_monitor_606);
    sample_manager_inst.add_one_monitor(fifo_monitor_607);
    sample_manager_inst.add_one_monitor(fifo_monitor_608);
    sample_manager_inst.add_one_monitor(fifo_monitor_609);
    sample_manager_inst.add_one_monitor(fifo_monitor_610);
    sample_manager_inst.add_one_monitor(fifo_monitor_611);
    sample_manager_inst.add_one_monitor(fifo_monitor_612);
    sample_manager_inst.add_one_monitor(fifo_monitor_613);
    sample_manager_inst.add_one_monitor(fifo_monitor_614);
    sample_manager_inst.add_one_monitor(fifo_monitor_615);
    sample_manager_inst.add_one_monitor(fifo_monitor_616);
    sample_manager_inst.add_one_monitor(fifo_monitor_617);
    sample_manager_inst.add_one_monitor(fifo_monitor_618);
    sample_manager_inst.add_one_monitor(fifo_monitor_619);
    sample_manager_inst.add_one_monitor(fifo_monitor_620);
    sample_manager_inst.add_one_monitor(fifo_monitor_621);
    sample_manager_inst.add_one_monitor(fifo_monitor_622);
    sample_manager_inst.add_one_monitor(fifo_monitor_623);
    sample_manager_inst.add_one_monitor(fifo_monitor_624);
    sample_manager_inst.add_one_monitor(fifo_monitor_625);
    sample_manager_inst.add_one_monitor(fifo_monitor_626);
    sample_manager_inst.add_one_monitor(fifo_monitor_627);
    sample_manager_inst.add_one_monitor(fifo_monitor_628);
    sample_manager_inst.add_one_monitor(fifo_monitor_629);
    sample_manager_inst.add_one_monitor(fifo_monitor_630);
    sample_manager_inst.add_one_monitor(fifo_monitor_631);
    sample_manager_inst.add_one_monitor(fifo_monitor_632);
    sample_manager_inst.add_one_monitor(fifo_monitor_633);
    sample_manager_inst.add_one_monitor(fifo_monitor_634);
    sample_manager_inst.add_one_monitor(fifo_monitor_635);
    sample_manager_inst.add_one_monitor(fifo_monitor_636);
    sample_manager_inst.add_one_monitor(fifo_monitor_637);
    sample_manager_inst.add_one_monitor(fifo_monitor_638);
    sample_manager_inst.add_one_monitor(fifo_monitor_639);
    sample_manager_inst.add_one_monitor(fifo_monitor_640);
    sample_manager_inst.add_one_monitor(fifo_monitor_641);
    sample_manager_inst.add_one_monitor(fifo_monitor_642);
    sample_manager_inst.add_one_monitor(fifo_monitor_643);
    sample_manager_inst.add_one_monitor(fifo_monitor_644);
    sample_manager_inst.add_one_monitor(fifo_monitor_645);
    sample_manager_inst.add_one_monitor(fifo_monitor_646);
    sample_manager_inst.add_one_monitor(fifo_monitor_647);
    sample_manager_inst.add_one_monitor(fifo_monitor_648);
    sample_manager_inst.add_one_monitor(fifo_monitor_649);
    sample_manager_inst.add_one_monitor(fifo_monitor_650);
    sample_manager_inst.add_one_monitor(fifo_monitor_651);
    sample_manager_inst.add_one_monitor(fifo_monitor_652);
    sample_manager_inst.add_one_monitor(fifo_monitor_653);
    sample_manager_inst.add_one_monitor(fifo_monitor_654);
    sample_manager_inst.add_one_monitor(fifo_monitor_655);
    sample_manager_inst.add_one_monitor(fifo_monitor_656);
    sample_manager_inst.add_one_monitor(fifo_monitor_657);
    sample_manager_inst.add_one_monitor(fifo_monitor_658);
    sample_manager_inst.add_one_monitor(fifo_monitor_659);
    sample_manager_inst.add_one_monitor(fifo_monitor_660);
    sample_manager_inst.add_one_monitor(fifo_monitor_661);
    sample_manager_inst.add_one_monitor(fifo_monitor_662);
    sample_manager_inst.add_one_monitor(fifo_monitor_663);
    sample_manager_inst.add_one_monitor(fifo_monitor_664);
    sample_manager_inst.add_one_monitor(fifo_monitor_665);
    sample_manager_inst.add_one_monitor(fifo_monitor_666);
    sample_manager_inst.add_one_monitor(fifo_monitor_667);
    sample_manager_inst.add_one_monitor(fifo_monitor_668);
    sample_manager_inst.add_one_monitor(fifo_monitor_669);
    sample_manager_inst.add_one_monitor(fifo_monitor_670);
    sample_manager_inst.add_one_monitor(fifo_monitor_671);
    sample_manager_inst.add_one_monitor(fifo_monitor_672);
    sample_manager_inst.add_one_monitor(fifo_monitor_673);
    sample_manager_inst.add_one_monitor(fifo_monitor_674);
    sample_manager_inst.add_one_monitor(fifo_monitor_675);
    sample_manager_inst.add_one_monitor(fifo_monitor_676);
    sample_manager_inst.add_one_monitor(fifo_monitor_677);
    sample_manager_inst.add_one_monitor(fifo_monitor_678);
    sample_manager_inst.add_one_monitor(fifo_monitor_679);
    sample_manager_inst.add_one_monitor(fifo_monitor_680);
    sample_manager_inst.add_one_monitor(fifo_monitor_681);
    sample_manager_inst.add_one_monitor(fifo_monitor_682);
    sample_manager_inst.add_one_monitor(fifo_monitor_683);
    sample_manager_inst.add_one_monitor(fifo_monitor_684);
    sample_manager_inst.add_one_monitor(fifo_monitor_685);
    sample_manager_inst.add_one_monitor(fifo_monitor_686);
    sample_manager_inst.add_one_monitor(fifo_monitor_687);
    sample_manager_inst.add_one_monitor(fifo_monitor_688);
    sample_manager_inst.add_one_monitor(fifo_monitor_689);
    sample_manager_inst.add_one_monitor(fifo_monitor_690);
    sample_manager_inst.add_one_monitor(fifo_monitor_691);
    sample_manager_inst.add_one_monitor(fifo_monitor_692);
    sample_manager_inst.add_one_monitor(fifo_monitor_693);
    sample_manager_inst.add_one_monitor(fifo_monitor_694);
    sample_manager_inst.add_one_monitor(fifo_monitor_695);
    sample_manager_inst.add_one_monitor(fifo_monitor_696);
    sample_manager_inst.add_one_monitor(fifo_monitor_697);
    sample_manager_inst.add_one_monitor(fifo_monitor_698);
    sample_manager_inst.add_one_monitor(fifo_monitor_699);
    sample_manager_inst.add_one_monitor(fifo_monitor_700);
    sample_manager_inst.add_one_monitor(fifo_monitor_701);
    sample_manager_inst.add_one_monitor(fifo_monitor_702);
    sample_manager_inst.add_one_monitor(fifo_monitor_703);
    sample_manager_inst.add_one_monitor(fifo_monitor_704);
    sample_manager_inst.add_one_monitor(fifo_monitor_705);
    sample_manager_inst.add_one_monitor(fifo_monitor_706);
    sample_manager_inst.add_one_monitor(fifo_monitor_707);
    sample_manager_inst.add_one_monitor(fifo_monitor_708);
    sample_manager_inst.add_one_monitor(fifo_monitor_709);
    sample_manager_inst.add_one_monitor(fifo_monitor_710);
    sample_manager_inst.add_one_monitor(fifo_monitor_711);
    sample_manager_inst.add_one_monitor(fifo_monitor_712);
    sample_manager_inst.add_one_monitor(fifo_monitor_713);
    sample_manager_inst.add_one_monitor(fifo_monitor_714);
    sample_manager_inst.add_one_monitor(fifo_monitor_715);
    sample_manager_inst.add_one_monitor(fifo_monitor_716);
    sample_manager_inst.add_one_monitor(fifo_monitor_717);
    sample_manager_inst.add_one_monitor(fifo_monitor_718);
    sample_manager_inst.add_one_monitor(fifo_monitor_719);
    sample_manager_inst.add_one_monitor(fifo_monitor_720);
    sample_manager_inst.add_one_monitor(fifo_monitor_721);
    sample_manager_inst.add_one_monitor(fifo_monitor_722);
    sample_manager_inst.add_one_monitor(fifo_monitor_723);
    sample_manager_inst.add_one_monitor(fifo_monitor_724);
    sample_manager_inst.add_one_monitor(fifo_monitor_725);
    sample_manager_inst.add_one_monitor(fifo_monitor_726);
    sample_manager_inst.add_one_monitor(fifo_monitor_727);
    sample_manager_inst.add_one_monitor(fifo_monitor_728);
    sample_manager_inst.add_one_monitor(fifo_monitor_729);
    sample_manager_inst.add_one_monitor(fifo_monitor_730);
    sample_manager_inst.add_one_monitor(fifo_monitor_731);
    sample_manager_inst.add_one_monitor(fifo_monitor_732);
    sample_manager_inst.add_one_monitor(fifo_monitor_733);
    sample_manager_inst.add_one_monitor(fifo_monitor_734);
    sample_manager_inst.add_one_monitor(fifo_monitor_735);
    sample_manager_inst.add_one_monitor(fifo_monitor_736);
    sample_manager_inst.add_one_monitor(fifo_monitor_737);
    sample_manager_inst.add_one_monitor(fifo_monitor_738);
    sample_manager_inst.add_one_monitor(fifo_monitor_739);
    sample_manager_inst.add_one_monitor(fifo_monitor_740);
    sample_manager_inst.add_one_monitor(fifo_monitor_741);
    sample_manager_inst.add_one_monitor(fifo_monitor_742);
    sample_manager_inst.add_one_monitor(fifo_monitor_743);
    sample_manager_inst.add_one_monitor(fifo_monitor_744);
    sample_manager_inst.add_one_monitor(fifo_monitor_745);
    sample_manager_inst.add_one_monitor(fifo_monitor_746);
    sample_manager_inst.add_one_monitor(fifo_monitor_747);
    sample_manager_inst.add_one_monitor(fifo_monitor_748);
    sample_manager_inst.add_one_monitor(fifo_monitor_749);
    sample_manager_inst.add_one_monitor(fifo_monitor_750);
    sample_manager_inst.add_one_monitor(fifo_monitor_751);
    sample_manager_inst.add_one_monitor(fifo_monitor_752);
    sample_manager_inst.add_one_monitor(fifo_monitor_753);
    sample_manager_inst.add_one_monitor(fifo_monitor_754);
    sample_manager_inst.add_one_monitor(fifo_monitor_755);
    sample_manager_inst.add_one_monitor(fifo_monitor_756);
    sample_manager_inst.add_one_monitor(fifo_monitor_757);
    sample_manager_inst.add_one_monitor(fifo_monitor_758);
    sample_manager_inst.add_one_monitor(fifo_monitor_759);
    sample_manager_inst.add_one_monitor(fifo_monitor_760);
    sample_manager_inst.add_one_monitor(fifo_monitor_761);
    sample_manager_inst.add_one_monitor(fifo_monitor_762);
    sample_manager_inst.add_one_monitor(fifo_monitor_763);
    sample_manager_inst.add_one_monitor(fifo_monitor_764);
    sample_manager_inst.add_one_monitor(fifo_monitor_765);
    sample_manager_inst.add_one_monitor(fifo_monitor_766);
    sample_manager_inst.add_one_monitor(fifo_monitor_767);
    sample_manager_inst.add_one_monitor(fifo_monitor_768);
    sample_manager_inst.add_one_monitor(fifo_monitor_769);
    sample_manager_inst.add_one_monitor(fifo_monitor_770);
    sample_manager_inst.add_one_monitor(fifo_monitor_771);
    sample_manager_inst.add_one_monitor(fifo_monitor_772);
    sample_manager_inst.add_one_monitor(fifo_monitor_773);
    sample_manager_inst.add_one_monitor(fifo_monitor_774);
    sample_manager_inst.add_one_monitor(fifo_monitor_775);
    sample_manager_inst.add_one_monitor(fifo_monitor_776);
    sample_manager_inst.add_one_monitor(fifo_monitor_777);
    sample_manager_inst.add_one_monitor(fifo_monitor_778);
    sample_manager_inst.add_one_monitor(fifo_monitor_779);
    sample_manager_inst.add_one_monitor(fifo_monitor_780);
    sample_manager_inst.add_one_monitor(fifo_monitor_781);
    sample_manager_inst.add_one_monitor(fifo_monitor_782);
    sample_manager_inst.add_one_monitor(fifo_monitor_783);
    sample_manager_inst.add_one_monitor(fifo_monitor_784);
    sample_manager_inst.add_one_monitor(fifo_monitor_785);
    sample_manager_inst.add_one_monitor(fifo_monitor_786);
    sample_manager_inst.add_one_monitor(fifo_monitor_787);
    sample_manager_inst.add_one_monitor(fifo_monitor_788);
    sample_manager_inst.add_one_monitor(fifo_monitor_789);
    sample_manager_inst.add_one_monitor(fifo_monitor_790);
    sample_manager_inst.add_one_monitor(fifo_monitor_791);
    sample_manager_inst.add_one_monitor(fifo_monitor_792);
    sample_manager_inst.add_one_monitor(fifo_monitor_793);
    sample_manager_inst.add_one_monitor(fifo_monitor_794);
    sample_manager_inst.add_one_monitor(fifo_monitor_795);
    sample_manager_inst.add_one_monitor(fifo_monitor_796);
    sample_manager_inst.add_one_monitor(fifo_monitor_797);
    sample_manager_inst.add_one_monitor(fifo_monitor_798);
    sample_manager_inst.add_one_monitor(fifo_monitor_799);
    sample_manager_inst.add_one_monitor(fifo_monitor_800);
    sample_manager_inst.add_one_monitor(fifo_monitor_801);
    sample_manager_inst.add_one_monitor(fifo_monitor_802);
    sample_manager_inst.add_one_monitor(fifo_monitor_803);
    sample_manager_inst.add_one_monitor(fifo_monitor_804);
    sample_manager_inst.add_one_monitor(fifo_monitor_805);
    sample_manager_inst.add_one_monitor(fifo_monitor_806);
    sample_manager_inst.add_one_monitor(fifo_monitor_807);
    sample_manager_inst.add_one_monitor(fifo_monitor_808);
    sample_manager_inst.add_one_monitor(fifo_monitor_809);
    sample_manager_inst.add_one_monitor(fifo_monitor_810);
    sample_manager_inst.add_one_monitor(fifo_monitor_811);
    sample_manager_inst.add_one_monitor(fifo_monitor_812);
    sample_manager_inst.add_one_monitor(fifo_monitor_813);
    sample_manager_inst.add_one_monitor(fifo_monitor_814);
    sample_manager_inst.add_one_monitor(fifo_monitor_815);
    sample_manager_inst.add_one_monitor(fifo_monitor_816);
    sample_manager_inst.add_one_monitor(fifo_monitor_817);
    sample_manager_inst.add_one_monitor(fifo_monitor_818);
    sample_manager_inst.add_one_monitor(fifo_monitor_819);
    sample_manager_inst.add_one_monitor(fifo_monitor_820);
    sample_manager_inst.add_one_monitor(fifo_monitor_821);
    sample_manager_inst.add_one_monitor(fifo_monitor_822);
    sample_manager_inst.add_one_monitor(fifo_monitor_823);
    sample_manager_inst.add_one_monitor(fifo_monitor_824);
    sample_manager_inst.add_one_monitor(fifo_monitor_825);
    sample_manager_inst.add_one_monitor(fifo_monitor_826);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(process_monitor_6);
    sample_manager_inst.add_one_monitor(process_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_8);
    sample_manager_inst.add_one_monitor(process_monitor_9);
    sample_manager_inst.add_one_monitor(process_monitor_10);
    sample_manager_inst.add_one_monitor(process_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
